���'     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.1�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i4�����R�(K�<�NNNJ����J����K t�b�C          �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h2�f8�����R�(KhKNNNJ����J����K t�b�C              �?       @�t�bhOh&�scalar���h2�i8�����R�(KhKNNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hK�
node_count�M��nodes�h(h+K ��h-��R�(KM���h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hhcK ��h�hcK��h�hcK��h�h[K��h�h[K ��h�hcK(��h�h[K0��uK8KKt�b�B�b         \                   @E@�J�+�?�           ��@       3                    �?+Jx��?L            @]@                           �?!Ce����?(             N@                          �_@hP�vCu�?            �D@                           �?�QN���?             ?@                           �?P���� �?             7@������������������������       �                      @       	                   �]@�G��l��?             5@������������������������       �                     @
                          `Z@��X��?	             ,@                          �Y@������?             @                          �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          ``@և���X�?             @                          �Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @                           �?���(\��?             $@                          �W@      �?             @������������������������       �                     �?                          �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          Pb@�q�q�?             @������������������������       �                     @������������������������       �                      @       $                   �Z@�p9W���?             3@        !                   �W@�8��8��?             @������������������������       �                     �?"       #                   @_@���Q��?             @������������������������       �                      @������������������������       �                     @%       .                   �`@8�Z$���?             *@&       +                    �?0�����?             @'       (                   0a@z�G�z�?             @������������������������       �                     @)       *                   `b@      �?              @������������������������       �                     �?������������������������       �                     �?,       -                    �?      �?              @������������������������       �                     �?������������������������       �                     �?/       2                   pb@      �?             @0       1                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @4       9                     �?���b���?$            �L@5       8                   @_@      �?             @6       7                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @:       ;                   �Z@�wN{/o�?             �J@������������������������       �                     ,@<       A                   �]@/y0��k�?            �C@=       >                   �]@؇���X�?             @������������������������       �                     @?       @                   �`@      �?             @������������������������       �                     �?������������������������       �                     @B       S                   �_@      �?             @@C       R                    �?��U�(�?             1@D       I                    \@�h$��W�?             .@E       H                    �?z�G�z�?             @F       G                   �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?J       Q                    @{�G�z�?             $@K       N                    ^@�n���?             "@L       M                   �`@VUUUUU�?             @������������������������       �      �?             @������������������������       �                      @O       P                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @T       [                    �?�r����?	             .@U       V                   0a@����X�?             @������������������������       �                     �?W       X                   �c@r�q��?             @������������������������       �                     @Y       Z                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @]       �                   �`@����V�?�           H�@^       g                   �U@h�T�B�?�            �n@_       f                    �?      �?              @`       a                   �a@�8��8��?             @������������������������       �                     @b       e                    �?�q�q�?             @c       d                   `e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @h       �                   �a@�M���?�            �m@i       z                     �?�Q����?d             d@j       s                    �?�q�����?             9@k       n                    _@�	j*D�?	             *@l       m                   Pr@      �?             @������������������������       �                     @������������������������       �                     �?o       r                    �?�����H�?             "@p       q                   `X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @t       u                    `@      �?	             (@������������������������       �                      @v       y                   �r@      �?             @w       x                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @{       �                   pa@l]?���?R            �`@|       �                   p`@6[�2���?B            @[@}       �                   �^@�R�Yߜ�?=            @Y@~                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �n@h�nOwA�?;            �X@�       �                    �?�~Q$�ɼ?'             Q@�       �                   �\@r�q��?             @������������������������       �                      @�       �                   pl@      �?             @�       �                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �h@���C�׷?#             O@�       �                    �?8�Z$���?             *@�       �                   @_@�8��8��?             (@������������������������       �                     "@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?@�E�x�?            �H@������������������������       �                     ?@�       �                    �?�X�<ݺ?             2@�       �                   �j@؇���X�?             @������������������������       �                      @�       �                    `@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                   �_@R���Q�?             >@�       �                   �n@�0�~�4�?             6@�       �                    �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     2@�       �                    �?      �?              @�       �                   �`@���Q��?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �b@      �?              @������������������������       �                     @�       �                    �?���Q��?             @�       �                    j@      �?             @������������������������       �                     �?�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?���B���?             :@�       �                   �e@     ��?
             0@������������������������       �                     @�       �                    �?���!pc�?             &@�       �                   �a@z�G�z�?             $@�       �                   �_@�<ݚ�?             "@������������������������       �                     @�       �                   0l@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?z�G�z�?             $@�       �                    ^@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �a@Hث3���?5            �S@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?�^B{	��?3             R@�       �                   �[@     ��?-             P@�       �                    X@ 	��p�?             =@������������������������       �                     *@�       �                   �e@      �?             0@������������������������       �                     �?�       �                    g@��S�ۿ?             .@������������������������       �        
             ,@������������������������       �                     �?�       �                   �\@���K�"�?            �A@�       �                    �?�$I�$I�?             @�       �                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    \@      �?             @�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?~h����?             <@�       �                    �?I�O���?             7@�       �                    �?�r����?             .@�       �                    h@r�q��?	             (@������������������������       �                      @������������������������       �                     $@������������������������       �                     @�       �                     �?      �?              @������������������������       �                      @�       �                   �e@�8��8��?             @�       �                   `b@      �?             @������������������������       �                     �?�       �                   0`@�q�q�?             @������������������������       �                     �?�       �                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @e@���Q��?             @�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    @      �?              @������������������������       �                     @�       �                     �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                  Pe@��� (�?�            0w@�       G                   �?�D���?�            0s@�       0                  Pc@JH�~�?N            ``@�       %                  0b@VUUUUe�?6             X@�                           �?��Ϙ#+�?-            @R@������������������������       �                     *@      $                  �b@�.�?��?&             N@      #                  8s@㜏u�?            �F@                        ``@���(\��?             D@                         ]@D'�$H{�?             =@                        �a@�z�G��?             $@                         �?      �?             @������������������������       �                      @                        �n@      �?             @	      
                  �m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @                         s@�*$�Z��?             3@                        �_@      �?
             0@                        �h@{�G�z�?             $@                        �_@      �?             @������������������������       �                     �?                        �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        a@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @                        �k@���!pc�?             &@                        �f@      �?             @������������������������       �                      @������������������������       �                      @                         �l@؇���X�?             @������������������������       �                     @!      "                  pa@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        	             .@&      '                  �b@Z��D�?	             7@������������������������       �                     @(      )                    �?��uJ���?             3@������������������������       �                     $@*      /                   �?VUUUUU�?             "@+      .                   �?      �?             @,      -                  �a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @1      F                  �r@E'���?            �A@2      =                  �`@n۶m۶�?             <@3      <                   _@     ��?             0@4      7                   �?      �?
             ,@5      6                  @]@z�G�z�?             @������������������������       �                     @������������������������       �                     �?8      ;                  e@�q�q�?             "@9      :                  �\@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @>      A                    �?      �?             (@?      @                   b@���Q��?             @������������������������       �                      @������������������������       �                     @B      C                  �i@����X�?             @������������������������       �                     �?D      E                  �c@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @H      k                  Pl@�X�B�?p             f@I      X                  �h@���F�?.            @Q@J      O                   �?�^�@�Y�?             =@K      N                   @      �?              @L      M                  �d@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @P      W                  `^@؇���X�?             5@Q      V                   @���Q��?             @R      S                   �?      �?             @������������������������       �                     �?T      U                  �g@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@Y      j                   �?      �?             D@Z      [                   �?�?�'�@�?             C@������������������������       �                     6@\      c                  �j@     ��?             0@]      b                  �j@և���X�?             @^      _                   @      �?             @������������������������       �                      @`      a                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @d      i                    �?�����H�?             "@e      h                  @_@z�G�z�?             @f      g                   k@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @l      �                   �?�3p�x��?B            �Z@m      ~                  �c@     ��?             @@n      {                  pc@�2'�%�?             7@o      r                   �?ƒ_,���?             .@p      q                  �b@      �?             @������������������������       �                     @������������������������       �                     �?s      v                  �_@���k���?             &@t      u                  8p@�q�q�?             @������������������������       �                     �?������������������������       �                      @w      z                   b@      �?              @x      y                  �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @|      }                   @      �?              @������������������������       �                     @������������������������       �                     �?      �                  �a@�����H�?             "@������������������������       �                      @������������������������       �                     �?�      �                   �?���9��?.            �R@�      �                  �b@أp=
��?(             N@�      �                  b@��S���?             .@�      �                   @���|���?	             &@�      �                  `]@�<ݚ�?             "@������������������������       �                     �?�      �                  �q@      �?              @������������������������       �                     @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                  �d@`Ӹ����?            �F@�      �                   @4?,R��?             B@�      �                  �c@     ��?             @@������������������������       �                     2@�      �                  �q@d}h���?
             ,@�      �                    �?և���X�?             @�      �                  �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   p@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                    �?      �?             @������������������������       �                      @������������������������       �                      @�      �                  0e@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�      �                  �_@���Q��?             .@������������������������       �                     @�      �                   b@"pc�
�?             &@�      �                  �o@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�      �                  �l@     �?(             P@�      �                  `f@      �?             @@������������������������       �        
             2@�      �                    @@4և���?             ,@������������������������       �                     *@������������������������       �                     �?�      �                  Pm@     `�?             @@������������������������       �                      @�      �                  `o@�h$���?             >@�      �                    �?B{	�%��?             "@������������������������       �                     @�      �                   �?      �?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  @_@      �?             @������������������������       �                      @�      �                  �`@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  �e@���N8�?             5@������������������������       �                     *@�      �                   �?      �?              @������������������������       �                     @�      �                  �q@      �?              @������������������������       �                     �?������������������������       �                     �?�t�b�values�h(h+K ��h-��R�(KM�KK��h[�BH*       �P@      x@     �q@      1@     �R@      :@      @     �A@      2@      @      <@      "@      @      8@      @      @      0@      @               @              @      ,@      @              @              @      @      @      @      @      �?              @      �?                      �?              @              @                              @      @              �?      @              �?                              @              @                       @              �?      @      @      �?       @      �?      �?                               @      �?                      �?               @                       @      @                      @               @              @      @      "@       @      @      �?                      �?       @      @               @                              @              �?      @       @      �?      �?      @              �?      @                      @              �?      �?              �?                              �?      �?              �?      �?                                      �?              @      @              @      �?                      �?              @                               @      $@     �C@       @      �?      �?       @      �?      �?                      �?              �?                                       @      "@      C@      @              ,@              "@      8@      @      @      �?              @                      @      �?                      �?              @                      @      7@      @      @      $@      @      @       @      @      �?      @              �?      @                      @              �?                              �?               @      @      @       @      @      @       @       @       @       @       @                               @              �?       @                       @              �?                      �?                       @                      *@       @              @       @                      �?              @      �?              @                      �?      �?                      �?              �?                       @             �H@     �s@      p@      8@     �f@      E@      @       @      @      �?       @      @                      @      �?       @              �?      �?              �?                              �?                      �?               @                      5@     @f@     �C@      "@     �_@      9@              (@      *@              "@      @              �?      @                      @              �?                       @      �?               @      �?                      �?               @                      @                      @      "@                       @              @      �?              �?      �?              �?                              �?               @              "@     �\@      (@      "@     @W@      @      "@      V@      @       @      �?                      �?               @                      @     �U@      @       @      P@       @      �?      @                       @              �?      @              �?      �?              �?                              �?                       @              �?     �M@       @              &@       @              &@      �?              "@                       @      �?                      �?               @                              �?      �?      H@                      ?@              �?      1@              �?      @                       @              �?      @              �?                              @                      &@              @      7@       @      �?      3@       @      �?      �?       @      �?      �?              �?                              �?                               @              2@              @      @               @      @               @       @                       @               @                              �?               @      �?                      �?               @                              @      @              @                       @      @               @       @              �?                      �?       @                       @              �?                              �?              5@      @              *@      @              @                       @      @               @       @              @       @              @                       @       @                       @               @                      �?                              �?               @       @              @       @              @                               @              @              (@      J@      ,@      @       @                       @              @                       @      I@      ,@      @     �H@      "@              ;@       @              *@                      ,@       @                      �?              ,@      �?              ,@                              �?      @      6@      @       @      �?      @      �?               @                       @      �?                      �?      �?       @      �?      �?              �?                              �?                               @      @      5@      @      @      2@      �?       @      *@               @      $@               @                              $@                      @               @      @      �?               @               @      @      �?       @       @                      �?               @      �?              �?                      �?      �?              �?                              �?                      �?      �?                      �?              �?                      @       @              �?       @              �?                               @               @               @      �?      @                      @       @      �?               @                              �?              9@     �`@     �j@      8@     �_@     �c@      *@     @S@     �D@      &@      O@      7@      @     �H@      4@              *@              @      B@      4@      @      5@      4@      @      0@      4@      @      *@      (@              @      @              @      @                       @              @      �?              �?      �?              �?                              �?               @                              @      @      $@      @      @      $@       @      @      @       @       @               @                      �?       @              �?                      �?       @                       @      @               @                              @                      @                              @              @       @               @       @                       @               @                      �?      @                      @              �?      @                      @              �?                      @                      .@              @      *@      @      @                      @      *@      @              $@              @      @      @              @      @              @      �?                      �?              @                               @      @                       @      .@      2@       @      .@      &@              @      "@              @      @              �?      @                      @              �?                      @      @              �?      @              �?                              @              @                               @       @       @       @       @      @               @                              @                      @       @                      �?              @      �?                      �?              @                              @      &@      I@     �\@      @      &@     �J@      @      @      2@      @      @              @      �?              @                              �?                       @                      @      2@              @       @              @      �?              �?                       @      �?               @                              �?                      �?                      0@              @     �A@              @     �@@                      6@              @      &@              @      @              �?      @                       @              �?      �?              �?                              �?              @                      �?       @              �?      @              �?      @                      @              �?                              �?                      @                       @      @     �C@      O@       @      1@      *@       @      "@      (@       @       @      @              �?      @                      @              �?               @      @       @       @              �?                      �?       @                              @      �?              �?      �?              �?                              �?              @                      �?      @                      @              �?                       @      �?               @                              �?      @      6@     �H@      @      *@     �E@               @      @              @      @               @      @              �?                      �?      @                      @              �?      �?                      �?              �?                       @                      @              @      @      B@              @      ?@              @      =@                      2@              @      &@              @      @               @      �?                      �?               @                      �?      @                      @              �?                              @               @       @                       @               @              @              @      @                                      @              "@      @                      @              "@       @              @       @              @                               @              @              �?      @      M@              �?      ?@                      2@              �?      *@                      *@              �?              �?      @      ;@               @              �?       @      ;@      �?      �?      @                      @      �?      �?      @              �?      �?              �?                              �?      �?              @                       @      �?              �?      �?                                      �?              �?      4@                      *@              �?      @                      @              �?      �?              �?                              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�Bg         j                   �^@�T!aA�?�           ��@       C                    `@��d���?V             a@                           Y@!���%�?)            @P@������������������������       �                      @       B                   �\@IӪ2�?%            �L@                           �?������?$            �K@������������������������       �                     @       !                    \@� 8o���?"            �I@	                           _@�8��8��?             8@
                          �Z@p=
ףp�?             $@                          `[@�8��8��?             @������������������������       �                      @                           �?      �?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                          �Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           D@������?	             ,@������������������������       �                      @                          b@�q�q�?             (@                           �?և���X�?             @                           �?z�G�z�?             @                          �W@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @                            �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @"       A                   @E@��1+��?             ;@#       $                   �Z@�+�wɃ�?             :@������������������������       �                     �?%       :                   �c@�^)��?             9@&       -                    �?b�2�tk�?             2@'       *                    ]@      �?             @(       )                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?+       ,                    _@      �?             @������������������������       �                     @������������������������       �                     �?.       9                   �^@�q�q�?             (@/       8                    �?      �?              @0       7                    �?և���X�?             @1       4                   `]@      �?             @2       3                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?5       6                     �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @;       >                    �?և���X�?             @<       =                   Pe@�q�q�?             @������������������������       �                     �?������������������������       �                      @?       @                   �_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @D       U                    �?�Ɖ�؇�?-            �Q@E       T                   �d@�`�7��?            �E@F       S                   Pd@l^Tv_�?            �D@G       L                    �?�p=
ף�?             D@H       I                   `]@�<ݚ�?             2@������������������������       �        	             $@J       K                    �?      �?              @������������������������       �                     @������������������������       �                     @M       R                   �`@���7�?             6@N       O                     �?�C��2(�?             &@������������������������       �                     �?P       Q                    `@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?������������������������       �                      @V       i                   a@�X�C�?             <@W       b                    ^@ףp=
��?             4@X       ]                    �?9��8���?             (@Y       Z                   �`@���Q��?             @������������������������       �                     �?[       \                   �W@      �?             @������������������������       �                     �?������������������������       �                     @^       a                   �]@և���X�?             @_       `                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @c       h                   �_@      �?              @d       e                    �?      �?             @������������������������       �                      @f       g                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @k                         �`@R����?s           ��@l       �                    �? ��՗��?�            �l@m       �                   p`@��<b�?h            �d@n       q                   �Y@L��t"�?d            �c@o       p                    �?      �?              @������������������������       �                     @������������������������       �                     @r       �                    �?��D�T.�?a            �b@s       x                   �U@�qk�M2�?I            �]@t       w                   `S@���Q��?             @u       v                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @y       |                     �?D�'��?F            @\@z       {                   `X@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@}       ~                   �W@�e }�r�??            @Y@������������������������       �                     $@       �                   �q@�$�-�?;            �V@�       �                    �?�p=
�#�?4             T@�       �                   @o@      �?             8@�       �                    Y@�	j*D�?             *@������������������������       �                      @�       �                   �_@"pc�
�?             &@������������������������       �                     @�       �                    _@���Q��?             @�       �                    `@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �p@�C��2(�?             &@������������������������       �                     @�       �                   @`@z�G�z�?             @������������������������       �                     �?�       �                   q@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �p@�$I�$I�?&             L@�       �                   �[@����m�?#            �J@�       �                   0a@���N8�?             5@�       �                   Pn@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             ,@�       �                   �[@     `�?             @@������������������������       �                     �?�       �                   �e@��e���?             ?@�       �                   �a@      �?             @������������������������       �                      @������������������������       �                      @�       �                    `@ ;����?             ;@�       �                   @c@�nkK�?             7@������������������������       �                     6@������������������������       �                     �?�       �                   @`@      �?             @������������������������       �                      @�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �_@VUUUUU�?             @������������������������       �                     �?�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�eP*L��?             &@�       �                   �Z@      �?              @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                      @�       �                    s@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �h@     `�?             @@�       �                   @\@      �?             @������������������������       �                     �?�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �U@�m۶m��?             <@�       �                    U@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    `@.n���?             9@�       �                   `\@ףp=
�?             4@������������������������       �                     $@�       �                   @_@z�G�z�?	             $@������������������������       �                     �?�       �                   Xq@�����H�?             "@������������������������       �                     @�       �                   `c@z�G�z�?             @������������������������       �                     �?�       �                   �]@      �?             @������������������������       �                     �?�       �                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �a@���Q��?             @������������������������       �                      @�       �                   t@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?և���X�?             @�       �                    j@      �?             @������������������������       �                      @�       �                   �^@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?     ��?.             P@�       �                   P`@h���h�?             �E@�       �                   @]@��Zy�?            �C@�       �                    �?�[��"e�?             2@�       �                    g@���Q��?             @�       �                   `c@      �?             @�       �                    X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?�؉�؉�?
             *@�       �                   �j@      �?             @������������������������       �                      @������������������������       �                      @�       �                     �?B{	�%��?             "@�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?؇���X�?             @�       �                   @e@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?؇���X�?             5@������������������������       �                     @�       �                   �a@@�0�!��?             1@�       �                    �?���!pc�?             &@������������������������       �                     @�       �                   �_@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�                         �i@>F?�!��?             5@�       �                     �?:/����?             @������������������������       �                     �?�                         �b@�8��8��?             @                          �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        
             ,@      �                  �w@./[-D��?�            w@      y                  �c@dO�%f�?�            �v@      r                  s@}A_��?r            �e@                         �?�h�Ai�?i            �c@	                        pl@g\�5�?             :@
                         �?j�V���?             &@                         @�$I�$I�?             @                          �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @                          �?�.�?��?             .@������������������������       �                      @                         �?�؉�؉�?	             *@                         �?      �?             (@                         `@      �?              @������������������������       �                     @                         b@      �?             @������������������������       �                     @������������������������       �                     �?                        �a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?      k                   �?H��gƴ�?W            �`@      Z                  hp@>��3p�?N            @^@       A                  pl@Zc1�Xu�?A            @Y@!      <                  �j@     ��?'             P@"      ;                  �j@ �o_��?             I@#      0                   �?��|�5��?            �G@$      -                   �?�q�q�?
             5@%      &                    �?�q�q�?             2@������������������������       �                      @'      (                  �[@      �?             0@������������������������       �                     @)      *                  `g@$�q-�?             *@������������������������       �                     $@+      ,                  �h@�q�q�?             @������������������������       �                     �?������������������������       �                      @.      /                   b@�q�q�?             @������������������������       �                     �?������������������������       �                      @1      :                  �b@8�Z$���?             :@2      9                   �?�8��8��?             8@3      4                  pa@�����H�?             2@������������������������       �                     �?5      6                   �?�IєX�?             1@������������������������       �                     @7      8                  @e@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     @������������������������       �                      @������������������������       �                     @=      @                   �?@4և���?
             ,@>      ?                  �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@B      W                   b@���L�?            �B@C      L                  �m@j���� �?             A@D      E                  `b@      �?             (@������������������������       �                     @F      K                  �b@      �?             @G      J                  ``@      �?             @H      I                  0m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @M      N                   Z@�GN�z�?             6@������������������������       �                      @O      V                  �a@R���Q�?             4@P      Q                  0a@�z�G��?             $@������������������������       �                     @R      S                  �n@և���X�?             @������������������������       �                     @T      U                  Hp@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@X      Y                  �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @[      j                   �?z�G�z�?             4@\      ]                  ``@�S����?             3@������������������������       �                     @^      _                   a@      �?             (@������������������������       �                     �?`      c                  @a@"pc�
�?             &@a      b                  �p@      �?              @������������������������       �                     �?������������������������       �                     �?d      e                    �?�����H�?             "@������������������������       �                     @f      i                  �q@r�q��?             @g      h                  @q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?l      m                  �^@�eP*L��?	             &@������������������������       �                     @n      q                   �?      �?              @o      p                  �j@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @s      x                   �?؇���X�?	             ,@t      u                  �t@$�q-�?             *@������������������������       �                     $@v      w                  �u@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?z      �                  `r@j��J�D�?g            �g@{      �                   �?�Pvv9��?R            �b@|      �                  j@�+78�/�?M            �a@}      �                  �h@̄���?            �D@~      �                   �?��ͦ-��?             ;@      �                  Pg@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  Pd@      �?             8@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?���7�?	             6@�      �                  �\@�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@������������������������       �                     @������������������������       �        
             ,@�      �                  @r@�cJ�͆�?6            �X@�      �                    �?��||��?5            @X@�      �                  �e@B{	�%��?             B@�      �                  �p@<�;��?             :@�      �                  `a@�HP��?
             9@�      �                   �?"pc�
�?             6@������������������������       �                     $@�      �                  0d@�q�q�?             (@������������������������       �                      @�      �                   �?z�G�z�?             $@������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                     @�      �                  �j@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�      �                  �a@���Q��?             $@������������������������       �                     @������������������������       �                     @�      �                  `l@���-�h�?'            �N@�      �                   k@@4և���?	             ,@�      �                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�      �                  �`@{���&�?            �G@�      �                  `d@D'�$H{�?             =@�      �                  �\@z�G�z�?             $@������������������������       �                     @�      �                  Pp@�q�q�?             @������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                  �d@R��Xp�?             3@������������������������       �                     @�      �                   �?{�G�z�?	             .@������������������������       �                      @�      �                  `e@g\�5�?             *@������������������������       �                     @�      �                  �n@���(\��?             $@������������������������       �                     @�      �                   �?      �?             @������������������������       �                     @�      �                  p@VUUUUU�?             @�      �                  �f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                  �q@�����H�?             2@������������������������       �        
             ,@�      �                  r@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�      �                    �?�eP*L��?             &@�      �                   �?      �?             @������������������������       �                      @������������������������       �                      @�      �                  pa@և���X�?             @�      �                   �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �                  u@�?�|�?            �B@������������������������       �                     @@�      �                   ]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                   c@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B(,       �M@     �u@     �t@      7@     �R@     �C@      2@      9@      6@               @              2@      1@      6@      2@      .@      6@      @                      ,@      .@      6@      "@      $@      @      �?      @       @      �?      @       @               @              �?      �?       @              �?      �?              �?                              �?      �?              �?      �?                                      �?              @               @      @      @               @               @      �?      @      @              @      @              �?      �?              �?      �?                                      �?      @                                       @      @      �?                      �?              @                      @      @      1@      @      @      0@              �?              @      @      0@      @      �?      (@      �?      �?      @              �?      �?                      �?              �?              �?              @                      @      �?                      @               @      @              @      @              @      @              @      �?              �?      �?                                      �?       @               @                       @       @                                      �?      �?                                      @              @      @              �?       @              �?                               @               @       @               @                               @                      �?               @              @     �H@      1@      �?     �A@      @      �?     �A@      @      �?     �A@      @              ,@      @              $@                      @      @              @                              @      �?      5@              �?      $@                      �?              �?      "@                      "@              �?                              &@                              �?                       @      @      ,@      $@      @      @      $@      @      @      @               @      @              �?                      �?      @              �?                              @      @      @              @      �?                      �?              @                               @                      �?      @              �?      @                       @              �?      �?              �?                              �?                      @               @              B@     �p@     0r@      9@     �c@     �F@      5@     @_@      3@      5@     �^@      .@              @      @              @                              @      5@     �]@      $@      1@      X@      @      @       @              �?       @                       @              �?                       @                      ,@     �W@      @              &@      �?                      �?              &@              ,@     �T@      @              $@              ,@     @R@      @      "@     �P@      @      @      3@      �?      @      "@               @                       @      "@                      @               @      @               @       @               @                               @                      �?                      $@      �?              @                      @      �?              �?                      @      �?                      �?              @              @      H@      @      @     �G@       @              4@      �?              @      �?                      �?              @                      ,@              @      ;@      �?      �?                      @      ;@      �?       @       @                       @               @                      �?      9@      �?      �?      6@                      6@              �?                              @      �?               @                      �?      �?                      �?              �?              �?      �?      �?              �?              �?              �?      �?                                      �?      @      @               @      @              �?                      �?      @                       @              �?      @                      @              �?                      @                      @      7@      @       @      �?      �?                      �?       @      �?                      �?               @                       @      6@      @              �?       @              �?                               @       @      5@       @              2@       @              $@                       @       @                      �?               @      �?              @                      @      �?              �?                      @      �?              �?                       @      �?                      �?               @               @      @                       @               @      �?               @                              �?                      @      @              @      @               @                      �?      @                      @              �?                              �?      @      A@      :@      �?      2@      8@      �?      ,@      8@      �?      &@      @               @      @               @       @              �?       @              �?                               @              �?                              �?      �?      "@      @               @       @               @                               @      �?      @      �?      �?      �?                      �?              �?                              @      �?              @      �?              @                              �?               @                      @      2@                      @              @      ,@              @       @                      @              @      @              @                              @                      @              @              @      0@       @      @       @       @              �?              @      �?       @      @      �?                      �?              @                                       @              ,@              &@      \@     �n@      &@     @Z@     �n@      @     �P@     @Y@      @     @P@     @V@       @      *@      &@      �?       @       @      �?      @       @      �?               @      �?                                       @              @                      @              �?      @      "@               @              �?      @      "@              @      "@              �?      @                      @              �?      @                      @              �?                       @       @                       @               @              �?                       @      J@     �S@       @      G@     @R@       @      >@     @Q@              .@     �H@              ,@      B@              &@      B@              @      ,@              @      (@               @                      @      (@              @                      �?      (@                      $@              �?       @              �?                               @              �?       @              �?                               @              @      6@               @      6@               @      0@              �?                      �?      0@                      @              �?      "@              �?                              "@                      @               @                      @                      �?      *@              �?      �?              �?                              �?                      (@       @      .@      4@              ,@      4@              "@      @              @                      @      @              �?      @              �?       @                       @              �?                              �?               @                      @      1@               @                      @      1@              @      @                      @              @      @                      @              @      �?              @                              �?                      $@       @      �?                      �?               @                              0@      @              0@      @              @                      "@      @                      �?              "@       @              �?      �?              �?                              �?               @      �?              @                      @      �?               @      �?               @                              �?              @                              �?              @      @                      @              @       @              @       @              @                               @              @                       @      (@              �?      (@                      $@              �?       @              �?                               @              �?              @      C@     �a@      @     �B@     �Z@      @      @@     @Y@      �?      @     �B@      �?      @      7@               @      �?                      �?               @              �?      �?      6@      �?              �?      �?                                      �?              �?      5@              �?      1@              �?                              1@                      @                      ,@      @      =@      P@      @      ;@      P@       @      &@      7@       @      @      3@       @      @      3@              @      2@                      $@              @       @               @                       @       @                      @               @      @                      @               @      �?               @                              �?       @              �?       @                                      �?              �?                      @      @              @                              @      @      0@     �D@              �?      *@              �?      @              �?                              @                      "@      @      .@      <@      @      *@      (@               @       @                      @               @      @                      @               @      �?               @                              �?      @      &@      @              @              @      @      @               @              @      @      @      @                      �?      @      @              @              �?      �?      @                      @      �?      �?      �?      �?              �?                      �?      �?                              �?                       @      0@                      ,@               @       @               @                               @               @                      @      @               @       @                       @               @                      @      @              @       @              @                               @                       @              �?      B@                      @@              �?      @              �?                              @              @       @                       @              @        �t�bub��!     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�f         v                  �c@��x<���?�           ��@       �                   �`@l�,M0�?u           ��@       �                    �?&�	-Z�?�            �t@                            �?ĊiӞ��?�            �m@                           �?l��[B��?             =@������������������������       �                     @                          �`@���Q��?             9@                          0r@X�<ݚ�?             2@	                           �?�q�q�?             .@
                           ]@�q�q�?             (@������������������������       �                     @                           _@      �?              @������������������������       �                     @                          �k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @                          @P@T�6|��?�             j@������������������������       �                      @       Y                   `_@T.�@���?�            �i@       6                   �[@BI-�܃�?.             O@       /                   �o@X��t��?             7@                          �Y@���[���?             2@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @       &                    �?�.�?��?             .@       !                   �X@      �?              @                            X@      �?             @������������������������       �                     �?������������������������       �                     @"       #                   �\@      �?             @������������������������       �                      @$       %                   �V@      �?              @������������������������       �                     �?������������������������       �                     �?'       .                    �?0�����?             @(       )                   �Z@      �?             @������������������������       �                      @*       -                   @[@      �?             @+       ,                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?0       1                    �?z�G�z�?             @������������������������       �                      @2       5                    �?�q�q�?             @3       4                    Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?7       R                    �?��#ۊ7�?            �C@8       O                    _@ʻ����?             A@9       N                   pl@      �?             @@:       =                    �?��s����?             5@;       <                   0i@      �?             @������������������������       �                     @������������������������       �                     �?>       A                   �Z@@�0�!��?             1@?       @                    Y@      �?              @������������������������       �                     �?������������������������       �                     �?B       M                   �U@�r����?	             .@C       L                   `]@r�q��?             (@D       K                   �_@�<ݚ�?             "@E       J                    \@      �?              @F       G                   `\@r�q��?             @������������������������       �                     @H       I                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        	             &@P       Q                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?S       V                    �?���Q��?             @T       U                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?W       X                   @Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @Z                          �b@��ӭ���?b             b@[       b                    �?����cU�?I            �[@\       a                   �[@�ӭ�a��?             2@]       `                   �[@{�G�z�?             @^       _                    Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        	             *@c       z                   a@<&����?<             W@d       e                   �X@X�����?             F@������������������������       �                      @f       u                   �`@�<ݚ�?             B@g       r                   �p@���B���?             :@h       i                   �]@�C��2(�?             6@������������������������       �                     *@j       k                    �?�<ݚ�?             "@������������������������       �                     @l       q                   `[@�q�q�?             @m       n                   �_@�q�q�?             @������������������������       �                     �?o       p                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @s       t                    �?      �?             @������������������������       �                     @������������������������       �                     �?v       y                    �?���Q��?             $@w       x                    `@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                      @{       |                    `@@��8��?             H@������������������������       �                     G@}       ~                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `d@�	U��6�?             A@�       �                    �?�eP*L��?             &@�       �                    �?����X�?             @������������������������       �                     �?�       �                   �N@�q�q�?             @�       �                   Pd@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    S@      �?             @�       �                   @d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �[@�l/���?             7@�       �                   �g@"pc�
�?	             &@�       �                   �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?      �?	             (@�       �                   �]@h/�����?             "@������������������������       �                     @�       �                   �e@z�G�z�?             @������������������������       �                     @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    m@VUUUUU�?             @������������������������       �                     �?�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��;�?=             W@�       �                   �X@     ��?             @@������������������������       �                     @�       �                    �?V�a�� �?             =@������������������������       �                     �?�       �                    �?�>4և��?             <@������������������������       �        
             0@�       �                   pa@�q�q�?             (@������������������������       �                     @�       �                   @^@      �?              @�       �                   8r@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �_@���ĳ��?)             N@�       �                    Z@���Er�?             1@������������������������       �                     �?�       �                   �U@     ��?             0@������������������������       �                      @�       �                   �o@d}h���?	             ,@�       �                     �?�8��8��?             (@������������������������       �                     @�       �                    \@�����H�?             "@�       �                   @\@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   @e@xa@��M�?            �E@�       �                    @      �?             E@�       �                    �?<�:�k+�?             ?@�       �                     �?�i�V��?             6@������������������������       �                     @�       �                    �?K&:~��?             3@�       �                   `c@�.�?��?             .@�       �                   s@r�q��?             (@�       �                    \@��!pc�?             &@������������������������       �                     �?�       �                   @_@ףp=
�?             $@������������������������       �                     @�       �                   @a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                    [@"pc�
�?             &@������������������������       �                      @�       �                   �a@�q�q�?             "@������������������������       �                     �?�       �                   �i@      �?              @�       �                    X@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       '                   �?ǵ@�A�?�            �m@�                          �a@�Yg}���?G            @\@�       �                    �?�������?             �I@�       �                    k@4��ݷ�?            �E@�       �                   �`@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                   �k@     `�?             @@������������������������       �                     @�       �                   �l@$I�$I��?             <@������������������������       �                     @�       �                   �`@      �?             8@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                     �?�&%�ݒ�?             5@������������������������       �                     @�       �                   �m@b�2�tk�?             2@������������������������       �                     @�       �                   @_@*D>��?
             *@�       �                    �?      �?              @�       �                   Hp@      �?             @�       �                   �o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �n@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �s@z�G�z�?             @������������������������       �                     @�       �                   �y@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �i@      �?              @������������������������       �                     @������������������������       �                     @                          �?�/�n�"�?'             O@                        0b@.k��\�?             1@������������������������       �                     @                         c@@4և���?
             ,@������������������������       �                     "@                        �q@z�G�z�?             @������������������������       �                      @                        pc@�q�q�?             @	      
                  0c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?      $                  Pc@X�<ݚ�?            �F@                         �?�q�q�?            �C@������������������������       �                     @                        0b@�<ݚ�?             B@                         �?�m۶m��?             <@                         �?j�V���?             6@                        �b@�lO���?             3@                        �a@�$I�$I�?             @������������������������       �                     @                        @_@      �?             @������������������������       �                     �?                        `g@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@                        `]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @       !                  �b@      �?              @������������������������       �                     @"      #                   �?���Q��?             @������������������������       �                      @������������������������       �                     @%      &                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @(      c                  pa@&3@�v��?R             _@)      0                  `Q@�`&�x��?7            �T@*      +                   �?      �?             @������������������������       �                     �?,      -                  �L@�q�q�?             @������������������������       �                     �?.      /                   �?      �?              @������������������������       �                     �?������������������������       �                     �?1      D                   �?vb'vb'�?3            �S@2      C                   �?l��\��?             A@3      4                  `a@�����H�?             ;@������������������������       �                     @5      6                   �?؇���X�?             5@������������������������       �                     �?7      B                   c@R���Q�?             4@8      A                  �p@z�G�z�?	             .@9      @                  b@؇���X�?             ,@:      ;                   l@      �?              @������������������������       �                     �?<      ?                  �a@؇���X�?             @=      >                  pn@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @E      L                   �?��ˠ�?             F@F      K                   �?p=
ףp�?             $@G      J                  �p@B{	�%��?             "@H      I                   \@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?M      T                  �j@�!���?             A@N      S                   �?�����H�?
             2@O      P                    �?"pc�
�?             &@������������������������       �                      @Q      R                  @e@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     @U      V                    �?     ��?             0@������������������������       �                      @W      b                   @X�Cc�?             ,@X      a                  �n@�eP*L��?	             &@Y      \                  `a@�q�q�?             "@Z      [                  �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @]      `                   b@r�q��?             @^      _                  l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @d      u                   �?�q�q�?             E@e      t                  xt@�z�G��?             D@f      s                  �q@�d�����?             C@g      l                   �?��}*_��?             ;@h      k                    �?�<ݚ�?             "@i      j                  �a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @m      n                   @r�q��?             2@������������������������       �                     (@o      r                   c@      �?             @p      q                  �]@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     &@������������������������       �                      @������������������������       �                      @w      �                   b@ħW1��?j             e@x      �                   @�:<����?Z            �a@y      �                  pl@*����?S            �`@z      �                    �?��4_O�?.            �S@{      �                  �a@      �?             8@|      }                   �?��Q��?             4@������������������������       �                     $@~                        @Y@�z�G��?             $@������������������������       �                      @�      �                   �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                  �P@�Jj�G�?!            �K@�      �                   �?��Q��?             $@������������������������       �                      @�      �                   �?      �?              @�      �                   �?������?             @�      �                  �[@�8��8��?             @������������������������       �                     @�      �                  Pe@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                   �?`Ӹ����?            �F@�      �                  �j@ףp=
�?             $@������������������������       �                     @�      �                   �?z�G�z�?             @������������������������       �                     @�      �                  ``@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  0d@��?^�k�?            �A@�      �                   �?�8��8��?             (@������������������������       �                     @�      �                  �j@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     7@�      �                   �?�1+�Q�?%             K@�      �                   �?���[���?             2@�      �                    �?ףp=
��?             $@�      �                  �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �d@և���X�?             @������������������������       �                     @�      �                  �p@      �?             @������������������������       �                     �?������������������������       �                     @�      �                   m@      �?              @������������������������       �                     �?�      �                  �\@؇���X�?             @������������������������       �                     @�      �                  @d@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   e@b�2�tk�?             B@�      �                  @_@��|���?             3@�      �                  �d@X�<ݚ�?             "@�      �                  pd@؇���X�?             @�      �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�      �                  d@z�G�z�?             $@������������������������       �                     @�      �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�      �                  �f@�t����?             1@������������������������       �        
             ,@�      �                  �s@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   a@�q�q�?             "@�      �                  �e@�q�q�?             @������������������������       �                     �?�      �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  `f@r�q��?             @�      �                  `a@�q�q�?             @������������������������       �                     �?�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                  �d@$�q-�?             :@������������������������       �                     6@�      �                  �e@      �?             @������������������������       �                      @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B�+       �H@     �v@      t@      C@     Pt@     `i@      <@      j@      W@      8@      e@     �F@              .@      ,@                      @              .@      $@               @      $@              @      $@              @      @              @                      �?      @                      @              �?       @              �?                               @                      @              @                      @              8@      c@      ?@                       @      8@      c@      =@      $@      C@      ,@      @      @      $@      @      @      $@               @      �?                      �?               @              @      �?      "@      @              @      @              �?                      �?      @                      �?              @                       @      �?              �?                      �?      �?                      �?      �?      @      �?      �?      @                       @      �?      �?       @      �?      �?              �?                              �?                               @                      �?      �?      @                       @              �?       @              �?      �?                      �?              �?                              �?              @      ?@      @      @      =@      �?      @      <@              @      1@              �?      @                      @              �?                      @      ,@              �?      �?                      �?              �?                       @      *@               @      $@               @      @              �?      @              �?      @                      @              �?       @              �?                               @                       @              �?                              @                      @                      &@                      �?      �?                      �?              �?                       @      @              �?      �?                      �?              �?                      �?       @              �?                               @      ,@     �\@      .@      @     �W@       @      �?      .@       @      �?       @       @      �?       @              �?                               @                               @              *@              @      T@      @      @     �@@      @               @              @      9@      @      @      5@               @      4@                      *@               @      @                      @               @      @               @      �?              �?                      �?      �?                      �?              �?                              @              @      �?              @                              �?                      @      @               @      @                      @               @                       @              �?     �G@                      G@              �?      �?                      �?              �?                      @      4@      @              @      @              @       @              �?                      @       @               @       @               @                               @               @                      �?      @              �?      �?                      �?              �?                               @      @      ,@       @       @      "@               @      �?                      �?               @                               @              @      @       @      @      @      �?      @                              @      �?              @                      �?      �?                      �?              �?              �?      �?      �?      �?                              �?      �?                      �?              �?              @     �D@     �G@              "@      7@              @                      @      7@              �?                      @      7@                      0@              @      @              @                      �?      @              �?      @              �?                              @                      @      @      @@      8@      �?      @      &@      �?                              @      &@               @                      @      &@              �?      &@                      @              �?       @              �?      @                       @              �?      �?                      �?              �?                              @               @              @      ;@      *@      @      ;@      (@      �?      5@      "@      �?      (@      "@              @              �?      "@      "@      �?      @      "@      �?       @      "@      �?      �?      "@              �?              �?              "@                      @      �?              @      �?                                      @              �?                      @                      @                      "@               @      @      @       @                              @      @                      �?              @       @               @       @               @                               @              @                              �?      $@      ]@     �[@      "@     @Q@     �A@      �?      :@      8@      �?      5@      5@              �?      $@              �?                              $@      �?      4@      &@              @              �?      0@      &@                      @      �?      0@      @              �?       @              �?                               @      �?      .@      @              @              �?      (@      @              @              �?      @      @              @      @              �?      @              �?      �?                      �?              �?                               @               @       @                       @               @              �?      @                      @              �?      �?              �?                              �?                      @      @              @                              @       @     �E@      &@      @      *@      �?      @                              *@      �?              "@                      @      �?               @                       @      �?              �?      �?              �?                              �?              �?              @      >@      $@      @      <@      @              @              @      9@      @       @      6@      @       @      0@      @      �?      0@       @      �?      @       @              @              �?      �?       @      �?                              �?       @                       @              �?                      (@              �?               @                       @      �?                              @              @      @       @      @                              @       @                       @              @                       @      @                      @               @              �?     �G@      S@      �?      3@      O@              @      �?              �?                       @      �?              �?                      �?      �?              �?                              �?      �?      0@     �N@              @      ?@              @      8@                      @              @      2@                      �?              @      1@              @      (@               @      (@               @      @              �?                      �?      @              �?      @                      @              �?                              @                      @              �?                              @                      @      �?      *@      >@      �?       @      @      �?      �?      @              �?      @              �?                              @      �?                              �?                      &@      7@               @      0@               @      "@                       @               @      @               @                              @                      @              "@      @                       @              "@      @              @      @              @      @              �?       @              �?                               @              @      �?               @      �?               @                              �?              @                               @              @                      <@      ,@              <@      (@              <@      $@              1@      $@               @      @               @       @                       @               @                              @              .@      @              (@                      @      @              �?      @              �?                              @               @                      &@                               @                       @      &@      D@     @]@      &@      C@     @W@      &@      @@     �V@      @      *@     �M@      @      @      *@              @      *@                      $@              @      @                       @              @      �?              @                              �?      @                      @      @      G@      @      @      @                       @      @      @      �?      @      @      �?      @       @      �?      @                               @      �?               @                              �?              �?                      �?                       @     �E@              �?      "@                      @              �?      @                      @              �?      �?              �?                              �?              �?      A@              �?      &@                      @              �?       @                       @              �?                              7@      @      3@      ?@       @      "@      @       @      @      @       @              �?                      �?       @                              @      @                      @              @      �?                      �?              @                      @       @                      �?              @      �?              @                       @      �?               @                              �?       @      $@      8@       @       @      "@       @      @      �?              @      �?               @      �?                      �?               @                      @               @                               @       @                      @               @      @               @                              @               @      .@                      ,@               @      �?                      �?               @                      @      @              �?       @                      �?              �?      �?                      �?              �?                      @      �?               @      �?              �?                      �?      �?                      �?              �?                      @                       @      8@                      6@               @       @               @                               @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�b         d                   �?�q���?�           ��@       =                   �c@�~�<��?u           ��@       (                    �?G��0��?4            @T@                          `]@,+}j��?&            �M@������������������������       �                     &@                            �?VUUUU��?             H@������������������������       �                     �?                          �_@��t2�?            �G@	                           I@��0f߻�?            �A@
                          �]@lxz�,C�?             9@                           �?     ��?             0@                          �[@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?������?
             ,@                           �?      �?              @                          p`@0�����?             @                          �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                          �W@VUUUUU�?             @������������������������       �                      @                          @`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@������������������������       �                     $@       %                   �`@      �?             (@       "                    �?������?             @        !                    d@      �?              @������������������������       �                     �?������������������������       �                     �?#       $                    �?���Q��?             @������������������������       �                      @������������������������       �                     @&       '                   �c@���Q��?             @������������������������       �                     @������������������������       �                      @)       4                    �?��!pc�?             6@*       -                   �]@{�G�z�?             .@+       ,                   @_@      �?              @������������������������       �                     �?������������������������       �                     @.       3                    �?և���X�?             @/       2                   `_@�q�q�?             @0       1                   P`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?5       <                   @e@և���X�?             @6       7                    `@z�G�z�?             @������������������������       �                      @8       ;                   `Q@�q�q�?             @9       :                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @>       �                     �?�6�i-�?A            ~@?       l                   �c@DA��ɒ�?U            ``@@       Q                    �?4.("�?9            @U@A       F                    _@\��"e��?             B@B       C                   �[@      �?             @������������������������       �                     �?D       E                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @G       N                   `c@     ��?             @@H       M                   �`@h�����?             <@I       J                    �?�����H�?             "@������������������������       �                      @K       L                   @Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             3@O       P                    �?      �?             @������������������������       �                     �?������������������������       �                     @R       g                    @և���X�?#            �H@S       T                   �g@�zv�X�?             F@������������������������       �                     @U       d                   hr@#z�i��?            �D@V       [                    �?�P�*�?             ?@W       X                   �\@     ��?	             0@������������������������       �                      @Y       Z                   �a@X�Cc�?             ,@������������������������       �                     "@������������������������       �                     @\       c                   Hq@��S���?             .@]       ^                   `i@�z�G��?	             $@������������������������       �                      @_       `                   �^@      �?              @������������������������       �                      @a       b                   �Z@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @e       f                    ^@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@h       k                    `@�Q����?             @i       j                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @m       �                   @|@v[X���?             G@n       y                   0e@
��N'�?            �F@o       x                   e@�ՙ/�?             5@p       s                    �?�"�O�|�?             1@q       r                   pd@�q�q�?             @������������������������       �                     �?������������������������       �                      @t       u                   �d@؇���X�?	             ,@������������������������       �                     &@v       w                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @z       {                    �? �q�q�?             8@������������������������       �        	             3@|       }                    ]@z�G�z�?             @������������������������       �                     �?~       �                    @      �?             @       �                   �e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       9                   �?d^o]�?�            �u@�       �                   �`@����w�?�             r@�       �                   hr@NW�0܋�?D            �Y@�       �                   �q@f?8���?9            �U@�       �                   �e@x����?7            �T@�       �                   �d@��(\�B�?5             T@�       �                    �?ʻ�
Wv�?4            �S@�       �                    c@�� �JH�?'            �M@�       �                    �?�3��?%            �L@�       �                   �Y@     ��?             0@������������������������       �                      @�       �                   p`@����S�?
             ,@�       �                   �k@�C��2(�?             &@������������������������       �                     @�       �                    _@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   @^@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   `_@̄���?            �D@�       �                   �k@�%d���?             =@�       �                   k@      �?             0@������������������������       �                     &@�       �                   �Y@�Q����?             @������������������������       �                     �?�       �                   0k@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             *@�       �                   �h@r�q��?             (@������������������������       �                      @������������������������       �                     $@�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��Q��?             4@�       �                   �m@      �?              @������������������������       �                     @�       �                   @[@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @`@�q�q�?	             (@�       �                   �`@�z�G��?             $@������������������������       �                     @�       �                   `b@      �?             @������������������������       �                      @�       �                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   (r@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     0@�                         e@$;=��?�             g@�                         �d@&���%(�?Y            �`@�       �                   �m@     b�?V             `@�       �                   pl@��"�O��?/             Q@�       �                    �?���QI�?&             I@�       �                   �[@���(\��?             4@�       �                   0j@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �_@���ĳ��?             .@�       �                   0a@:/����?             @������������������������       �                     �?�       �                   �a@�8��8��?             @�       �                   �a@      �?             @�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   0k@      �?              @�       �                   0c@؇���X�?             @�       �                    b@�q�q�?             @������������������������       �                     �?�       �                   `g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �a@z�G�z�?             >@������������������������       �                     *@�       �                   �k@ҳ�wY;�?             1@�       �                    �?և���X�?             ,@������������������������       �                      @�       �                   @e@�q�q�?             (@������������������������       �                     �?�       �                   �_@���!pc�?
             &@�       �                   c@      �?             @�       �                   �\@���Q��?             @������������������������       �                     �?�       �                   b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?&���^B�?	             2@�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   m@      �?             0@�       �                   �l@���Q��?             $@������������������������       �                     @�       �                    ]@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�                         Pc@��A���?'             N@�                          �?�"e����?             B@�       �                   �n@���[���?
             2@������������������������       �                      @�       �                   �o@     ��?	             0@������������������������       �                     @�                          �a@�	j*D�?             *@�       �                   �_@      �?             @������������������������       �                     @������������������������       �                     �?                        @^@�����H�?             "@                        �[@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                        �q@�<ݚ�?             2@                         \@      �?
             0@������������������������       �                     �?	                         �?��S�ۿ?	             .@
                        @`@      �?             @������������������������       �                      @                        b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                      @                         _@�8��8��?             8@                         �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     1@������������������������       �                     @                          �?�R�k���?(            �I@                        �f@�}�+r��?             3@                        Pf@؇���X�?             @������������������������       �                     @                         �?�q�q�?             @                        @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@!      6                   @      �?             @@"      %                  `]@H�7�&��?             >@#      $                  `\@      �?             @������������������������       �                     �?������������������������       �                     @&      +                   �?�K8��?             :@'      *                  (r@r�q��?             @(      )                  �o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @,      5                  �`@ףp=
�?             4@-      4                  @g@z�G�z�?
             $@.      3                   �?�����H�?	             "@/      2                  @^@r�q��?             @0      1                  0e@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     $@7      8                  @`@      �?              @������������������������       �                     �?������������������������       �                     �?:      I                   `@$E��b��?'            �N@;      <                  @j@��e���?             ?@������������������������       �                     @=      H                  @^@�q�q�?             8@>      C                  Pm@.k��\�?             1@?      @                  �\@      �?             @������������������������       �                      @A      B                  �k@      �?              @������������������������       �                     �?������������������������       �                     �?D      E                  @e@$�q-�?             *@������������������������       �                     &@F      G                  �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @J      U                   �?d��0u��?             >@K      T                   a@�n_Y�K�?             *@L      M                  �`@X�<ݚ�?             "@������������������������       �                     �?N      O                  pa@      �?              @������������������������       �                     �?P      Q                  �m@և���X�?             @������������������������       �                      @R      S                  �n@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @V      ]                  ``@@�0�!��?             1@W      X                   �?����X�?             @������������������������       �                     @Y      Z                  `^@�q�q�?             @������������������������       �                     �?[      \                  Pb@      �?              @������������������������       �                     �?������������������������       �                     �?^      _                  @a@ףp=
�?             $@������������������������       �                     @`      c                   �?z�G�z�?             @a      b                  �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @e      �                  `_@��/��g�?j            �e@f      o                  �Y@lK���?             G@g      j                  `X@      �?              @h      i                  �`@      �?             @������������������������       �                     �?������������������������       �                     @k      n                   �?      �?             @l      m                  �\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?p      �                   �?��k(��?             C@q      t                    �?�'��P��?             ;@r      s                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @u      x                   \@e�J��?             5@v      w                  �Z@      �?             @������������������������       �                      @������������������������       �                      @y      z                  �Z@f�t���?             1@������������������������       �                     @{      |                  �]@�$I�$I�?	             ,@������������������������       �                     @}      �                  �^@��!pc�?             &@~                        �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �a@      �?              @������������������������       �                     @�      �                  Pe@      �?             @������������������������       �                     @������������������������       �                     �?�      �                   �?"pc�
�?             &@�      �                   e@z�G�z�?             $@�      �                   \@�q�q�?             @������������������������       �                     �?�      �                  �^@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   g@R�
S�{�?L            �_@�      �                  �d@�>��V�?K            @_@�      �                  �p@Z�����?B            @[@�      �                   �?�����?1            �T@�      �                   d@�J�4�?             I@�      �                   �?��S�ۿ?            �F@�      �                  @^@Pa�	�?            �@@������������������������       �        	             0@�      �                  �N@�IєX�?	             1@�      �                  c@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@�      �                  0i@r�q��?	             (@������������������������       �                     @�      �                   a@����X�?             @�      �                  Pb@���Q��?             @�      �                   �?      �?             @�      �                  �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                  @a@�U�I��?            �@@������������������������       �                     *@�      �                  �i@z�G�z�?             4@�      �                   �?>;n,��?             &@������������������������       �                     @�      �                  `a@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�      �                   �?��WV��?             :@�      �                   �?�S����?             3@�      �                  �]@�n���?             "@�      �                  @s@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                  �`@      �?             @�      �                  `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�      �                  `c@����X�?             @�      �                  �q@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �        	             0@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KM�KK��h[�BH*       �I@     0x@     �r@      >@     0q@      p@      &@      J@      2@      @      E@      $@              &@              @      ?@      $@                      �?      @      ?@      "@      @      <@      @      @      2@      @      @      "@      @      �?      �?              �?                              �?              @       @      @      �?      @      �?      �?      @      �?      �?              �?      �?                                      �?              @                      �?               @       @       @               @               @               @       @                                       @              "@                      $@              @      @      @      @      �?      @              �?      �?              �?                              �?      @               @                       @      @                               @      @                      @               @              @      $@       @      @      @      @      �?      @              �?                              @              @              @       @              @       @              @       @                                      @                      �?      �?                              @      @              �?      @                       @              �?       @              �?      �?              �?                              �?                      �?               @              3@     �k@     �m@      @      M@     �Q@       @      I@     �@@      �?      @@      @               @       @              �?                      �?       @              �?                               @      �?      >@      �?              ;@      �?               @      �?               @                      @      �?                      �?              @                      3@              �?      @              �?                              @              �?      2@      >@              1@      ;@              @                      ,@      ;@              *@      2@              @      &@                       @              @      "@                      "@              @                       @      @              @      @                       @              @      @               @                      �?      @              �?                              @              @                      �?      "@              �?                              "@      �?      �?      @      �?      �?                      �?              �?                                      @      �?       @     �B@      �?      @     �B@      �?      @      ,@      �?       @      ,@      �?               @      �?                                       @               @      (@                      &@               @      �?                      �?               @                      @                      �?      7@                      3@              �?      @                      �?              �?      @              �?       @                       @              �?                              �?              �?              0@     �d@      e@      .@     �_@     @b@       @     @R@      6@       @     �L@      6@      @     �L@      4@      @     �L@      1@      @     �L@      1@      @      I@      @      @     �H@      @      @      (@      �?       @                      �?      (@      �?      �?      $@                      @              �?      @              �?                              @                       @      �?                      �?               @              �?     �B@      @      �?      ;@      �?      �?      ,@      �?              &@              �?      @      �?                      �?      �?      @              �?                              @                      *@                      $@       @                       @              $@              �?      �?                      �?              �?                              @      *@               @      @                      @               @      �?               @                              �?              @      @              @      @                      @              @      �?               @                      �?      �?                      �?              �?                       @              �?                                      @       @               @       @                                       @              0@              @      K@      _@      @      H@     @T@      @      E@     @T@      @      ;@      C@       @      ,@      A@       @       @      $@              @      �?              @                              �?       @      @      "@       @       @      @      �?                      �?       @      @              �?      @              �?       @                       @              �?                              �?      �?      �?              �?                              �?                       @      @              �?      @              �?       @                      �?              �?      �?                      �?              �?                              @              �?                      @      8@                      *@              @      &@              @       @               @                      @       @              �?                      @       @              @      @               @      @                      �?               @       @               @                               @              �?                              @                      @      �?      *@      @      �?      �?              �?                              �?                      (@      @              @      @              @                       @      @               @                              @              @               @      .@     �E@       @      *@      5@       @      "@      @       @                              "@      @                      @              "@      @              �?      @                      @              �?                       @      �?              @      �?              @                              �?              @                      @      ,@               @      ,@              �?                      �?      ,@              �?      @                       @              �?      �?                      �?              �?                              &@               @                       @      6@               @      @               @                              @                      1@              @               @      @     �E@              �?      2@              �?      @                      @              �?       @              �?      �?                      �?              �?                              �?                      (@       @      @      9@       @      @      8@              @      �?                      �?              @               @      �?      7@              �?      @              �?       @                       @              �?                              @       @              2@       @               @      �?               @      �?              @      �?              @      �?                                      @                      �?                      @      �?                                      $@              �?      �?              �?                              �?      �?      C@      6@      �?      ;@      @              @              �?      4@      @      �?      *@      @      �?      �?       @                       @      �?      �?                      �?              �?                              (@      �?              &@                      �?      �?                      �?              �?                      @                      &@      3@               @      @              @      @              �?                      @      @                      �?              @      @               @                      �?      @                      @              �?                      @                      @      ,@               @      @                      @               @      �?              �?                      �?      �?              �?                              �?              �?      "@                      @              �?      @              �?       @                       @              �?                               @      5@      \@      D@      $@      *@      7@      @      @              @      �?                      �?              @                      �?      @              �?       @                       @              �?                              �?              @      "@      7@      @      @      ,@       @              @                      @       @                      @      @      $@       @               @                       @       @                       @      @       @              @               @      @       @                      @       @      @      @       @      �?                      �?               @                              @      @                      @              @      �?              @                              �?               @      "@               @       @               @      @              �?                      �?      @                      @              �?                              @                      �?      &@     �X@      1@      "@     �X@      1@      "@     �T@      1@      @     @Q@      "@              E@       @              E@      @              @@      �?              0@                      0@      �?              @      �?              @                              �?              &@                      $@       @              @                      @       @              @       @              @      �?               @      �?                      �?               @                      �?                              �?               @                              @      @      ;@      �?              *@              @      ,@      �?      @      @      �?              @              @              �?      @                                      �?              "@              @      ,@       @      @      (@      @      @       @      @      @      �?                      �?              @                              �?      @              �?      �?              �?                              �?                       @              $@                       @      @              �?      @              �?                              @              �?                      0@               @                �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�BXa         >                  c@�	v��?�           ��@                          `_@�*b7�U�?T           H�@       R                    �?g*�h�?q            @f@       C                    �?�{�yX�?K            �]@       *                   p`@�;fq��?;            �V@                           [@��e�S�?'            �L@                           �?&�q-�?             *@                           �?      �?              @	       
                   @l@      �?              @������������������������       �                     �?������������������������       �                     �?                          �\@�q�q�?             @������������������������       �                      @                          �Y@      �?             @������������������������       �                      @������������������������       �                      @                           �?�Q����?             @������������������������       �                     �?                          �Z@      �?             @������������������������       �                     @������������������������       �                     �?                           �?��Z=;�?             F@                          �R@@4և���?             <@                          �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     9@       )                   `]@     ��?
             0@       $                   `Z@�؉�؉�?             *@       !                    ]@{�G�z�?             @                           `[@      �?              @������������������������       �                     �?������������������������       �                     �?"       #                   `X@�q�q�?             @������������������������       �                     �?������������������������       �                      @%       (                   p`@      �?              @&       '                    \@z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �                     @+       B                   pb@&5DS�?             A@,       /                     �?��y�):�?             9@-       .                    Y@      �?             @������������������������       �                     @������������������������       �                     �?0       A                    b@�ՙ/�?             5@1       @                    �?X�<ݚ�?             2@2       3                   �`@j���� �?             1@������������������������       �                     �?4       5                    a@     ��?
             0@������������������������       �                     �?6       ;                   �o@���Q��?	             .@7       8                   �[@z�G�z�?             $@������������������������       �                     �?9       :                   �^@�����H�?             "@������������������������       �                      @������������������������       �                     �?<       ?                   �a@z�G�z�?             @=       >                   �p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@D       G                     �?�5��?             ;@E       F                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?H       Q                   @^@      �?             8@I       P                   �`@�GN��?             6@J       O                   8t@0�����?	             2@K       L                    X@�IєX�?             1@������������������������       �                      @M       N                   �\@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @S       `                    �?���(\��?&             N@T       Y                   `]@:/����?	             ,@U       V                     �?      �?             @������������������������       �                     �?W       X                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?Z       [                    ^@H�z�G�?             $@������������������������       �                     @\       _                   �^@������?             @]       ^                   �[@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @a       f                     �?
;&����?             G@b       c                   q@�t����?
             1@������������������������       �                     *@d       e                   q@      �?             @������������������������       �                      @������������������������       �                      @g       l                    \@Y��sd�?             =@h       i                   �X@      �?              @������������������������       �                     �?j       k                   �S@և���X�?             @������������������������       �                     @������������������������       �                     @m       ~                   �^@և���X�?             5@n       }                    @�\��N��?             3@o       v                   pk@     ��?             0@p       q                   �]@����X�?             @������������������������       �                     �?r       u                    �?r�q��?             @s       t                   �h@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @w       |                   �p@�<ݚ�?             "@x       y                    �?      �?              @������������������������       �                     @z       {                   �\@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?p����?�            pu@�       �                     �?�r)��?�            �l@�       �                    �?      �?             @@������������������������       �                      @�       �                   �m@ �q�q�?             8@�       �                    �?�8��8��?             (@�       �                   �`@ףp=
�?             $@�       �                   0k@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     (@�       �                   `@��aK]��?~            �h@�       �                    �?��3�͸�?U             `@�       �                    �?�����?;            �T@�       �                   �`@��e���?)             O@������������������������       �        
             .@�       �                   �`@�6f�+��?            �G@������������������������       �                     �?�       �                    �?Ļ��|�?             G@�       �                   �[@      �?             @������������������������       �                     �?�       �                    c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   0k@�p=
ף�?             D@�       �                   pe@/����?
             ,@������������������������       �                     $@�       �                   �]@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   0c@ ��WV�?             :@������������������������       �                     *@�       �                   �Z@$�q-�?             *@������������������������       �                     $@�       �                   Pd@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @R@>F?�!��?             5@������������������������       �                      @�       �                    ^@�lO���?             3@�       �                   �q@�8��8��?             (@������������������������       �        
             &@������������������������       �                     �?�       �                   `Y@����X�?             @�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �n@z�G�z�?             @������������������������       �                     @�       �                   `_@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   hq@��<b���?             G@�       �                    �?r�q��?             B@�       �                   �b@�z�G��?
             4@�       �                   �`@$�q-�?             *@�       �                    j@r�q��?             @������������������������       �                     @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �c@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@�       �                   �q@���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                    �? ���ٻ�?)            �P@�       �                    �?¦�F0�?            �D@�       �                   �j@"��u���?             9@�       �                   �`@      �?              @������������������������       �                     �?�       �                   Pi@؇���X�?             @�       �                    a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   0b@ҳ�wY;�?             1@�       �                   �r@؇���X�?             ,@������������������������       �                     "@�       �                   8s@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   Pm@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @d@     ��?	             0@�       �                   �`@�	j*D�?             *@������������������������       �                      @�       �                    g@"pc�
�?             &@������������������������       �                     @�       �                   �a@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �i@�n_Y�K�?             :@�       �                    �?��S�ۿ?             .@������������������������       �                     @�       �                   @W@�C��2(�?             &@�       �                    `@؇���X�?             @������������������������       �                     @�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   ``@�C��2(�?             &@�       �                   `c@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�                           �?�AbL���?Q            �\@�                           @(ݾ�z��?             :@�       �                   �\@8����?             7@������������������������       �                     @�       �                    a@z�G�z�?             4@������������������������       �                     "@�       �                   0a@���|���?             &@������������������������       �                     @�       �                   �s@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                         b@�q�q�?             @������������������������       �                     �?                        `c@      �?              @������������������������       �                     �?������������������������       �                     �?                         �?1T)�q�?>            @V@                         �?j�Y�H��?             >@      	                  �X@�;�;�?             :@������������������������       �                     �?
                        �`@`�Q��?             9@                        �`@B{	�%��?             "@                        ``@      �?              @                         W@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                        �n@      �?             0@������������������������       �        	             *@                        `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        �`@      �?             @������������������������       �                      @                         b@      �?              @������������������������       �                     �?������������������������       �                     �?      +                  P`@Z�ï:2�?%            �M@                        �V@.n���?             9@������������������������       �                     @      *                  �b@���(\��?	             4@       !                   `@X�<ݚ�?             2@������������������������       �                     �?"      )                  �a@j���� �?             1@#      $                  pm@�q�q�?             (@������������������������       �                      @%      (                  �`@�z�G��?             $@&      '                  �r@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @,      -                  0a@�"�O�|�?             A@������������������������       �        	             (@.      3                  �a@j�V���?             6@/      2                  �a@{�G�z�?             @0      1                  �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @4      =                  �^@@�0�!��?             1@5      6                   �?�θ�?	             *@������������������������       �                      @7      <                   �?���!pc�?             &@8      ;                  �j@�q�q�?             "@9      :                  `T@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @?      �                  �w@�lo���?�            �j@@      Q                  �c@H�K��%�?�             j@A      B                   �?�n_Y�K�?             *@������������������������       �                     �?C      P                   b@�q�q�?             (@D      O                  �Q@���!pc�?
             &@E      H                   �?�q�q�?             "@F      G                   e@      �?              @������������������������       �                     �?������������������������       �                     �?I      N                   �?����X�?             @J      K                  pc@      �?             @������������������������       �                     �?L      M                  �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?R      �                   @��G���?�            �h@S      �                   �?)�ݧ��?x            `g@T      �                  `f@�����8�?o            `e@U      �                  0e@�w��s��?l            �d@V      w                    �?�T���N�?C             Y@W      n                   �?��]�"�?            �C@X      m                  e@Hm���?             =@Y      b                   �?��P��?             ;@Z      a                   �?ףp=
��?             $@[      \                  `a@�8��8��?             @������������������������       �                      @]      ^                  �c@      �?             @������������������������       �                     �?_      `                  d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @c      f                   �?������?
             1@d      e                  �b@      �?             @������������������������       �                      @������������������������       �                      @g      h                  p@8�Z$���?             *@������������������������       �                      @i      j                  @`@���Q��?             @������������������������       �                      @k      l                  `b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @o      r                  @^@H�z�G�?             $@p      q                  �c@      �?             @������������������������       �                     @������������������������       �                     �?s      v                  Pd@r�q��?             @t      u                  �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @x      �                  �q@4-7nN,�?-            �N@y      �                  �d@���Er�?'            �I@z      {                  pi@�q�q�?              E@������������������������       �                      @|      �                  d@j���� �?             A@}      �                   �?�q�q�?             8@~      �                   �?�z�G��?             4@      �                  �c@����X�?             @������������������������       �                     @������������������������       �                      @�      �                  �p@�	j*D�?             *@������������������������       �                      @�      �                  �\@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                  �^@      �?             @������������������������       �                      @������������������������       �                      @�      �                  �k@���Q��?             $@������������������������       �                     @�      �                   �?؇���X�?             @�      �                   �?r�q��?             @�      �                  �o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                  @l@x�5?,�?             "@�      �                   �?      �?             @������������������������       �                      @�      �                  Pk@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  �o@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@�      �                   �?      �?)             P@�      �                  �q@     ��?             0@������������������������       �                     "@�      �                   f@����X�?             @�      �                  �r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                  �e@      �?             H@������������������������       �                     0@�      �                  @^@     ��?             @@�      �                    �?      �?	             (@�      �                  �i@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?z�G�z�?             $@������������������������       �                     @�      �                  `\@      �?             @�      �                  �f@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@������������������������       �                     @������������������������       �        	             0@�      �                  �j@�q�q�?             "@������������������������       �                      @�      �                  d@؇���X�?             @������������������������       �                     @�      �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B�)        K@     �v@     �s@      H@     @s@     �d@      8@     @T@     @R@      ,@     @P@     �C@      (@      M@      5@      "@     �D@      @      @      @      �?      @      @              �?      �?                      �?              �?                      @       @               @                       @       @                       @               @                      �?      @      �?                      �?      �?      @                      @              �?                      @     �A@      @              :@       @              �?       @              �?                               @              9@              @      "@      @      @      "@      �?       @       @      �?              �?      �?              �?                              �?       @      �?                      �?               @                      �?      @              �?      @                       @              �?       @                      @                              @      @      1@      ,@      @       @      ,@      @              �?      @                                      �?               @      *@               @      $@              @      $@                      �?              @      "@              �?                      @      "@               @       @              �?                      �?       @                       @              �?                      @      �?               @      �?               @                              �?               @                      �?                              @              "@               @      @      2@      �?               @                       @      �?                      �?      @      0@      �?      @      0@      �?      �?      0@      �?              0@                       @      �?               @                       @      �?                              �?                      @                       @              $@      0@      A@      @      @      @              @      �?              �?                       @      �?               @                              �?      @      �?      @      @                      @      �?      @              �?      @              �?                              @      @                      @      (@      >@               @      .@                      *@               @       @               @                               @      @      $@      .@      @      �?      @              �?              @              @      @                                      @              "@      (@              "@      $@              "@      @               @      @              �?                      �?      @              �?      �?              �?                              �?                      @              @       @              @      �?              @                      @      �?                      �?              @                              �?                      @                       @      8@     `l@      W@      2@     �e@     �B@              ?@      �?               @                      7@      �?              &@      �?              "@      �?              @      �?              @                              �?              @                       @                      (@              2@     �a@      B@      "@     �Z@      ,@      "@     �Q@      @      @      K@       @              .@              @     �C@       @      �?                      @     �C@       @      �?      @      �?                      �?      �?      @                      @              �?                      @     �A@      �?      @      $@      �?              $@              @              �?      @                                      �?      �?      9@                      *@              �?      (@                      $@              �?       @              �?                               @              @      0@       @       @                      �?      0@       @      �?      &@                      &@              �?                              @       @              �?      �?                      �?              �?                      @      �?              @                      �?      �?                      �?              �?                      B@      $@              >@      @              ,@      @              (@      �?              @      �?              @                       @      �?                      �?               @                      @                       @      @                      @               @                      0@                      @      @                      @              @              "@      B@      6@      @      2@      2@       @      ,@      "@               @      @              �?                      �?      @              �?       @                       @              �?                              @       @      (@      @              (@       @              "@                      @       @                       @              @               @              �?                      �?       @                      @      @      "@              @      "@               @                       @      "@                      @               @      @               @                              @      @                      @      2@      @      �?      ,@                      @              �?      $@              �?      @                      @              �?      @              �?                              @                      @              @      @      @      @      @              @                              @                      �?      @              �?      �?                      �?              �?                              @      @      K@     �K@      �?      @      2@              @      0@              @                      @      0@                      "@              @      @                      @              @      �?              @                              �?      �?               @                      �?      �?              �?      �?                                      �?      @     �G@     �B@      �?      @      7@      �?      @      6@              �?              �?       @      6@      �?      �?      @      �?              @      �?              @      �?                                      @                      �?              �?                      �?      .@                      *@              �?       @                       @              �?                      @      �?               @                      �?      �?                      �?              �?              @     �D@      ,@       @      *@      $@              @               @       @      $@               @      $@              �?                      @      $@              @      @                       @              @      @              �?      @                      @              �?                      @                              @       @                       @      <@      @              (@               @      0@      @       @       @      �?               @      �?                      �?               @               @                              ,@      @              $@      @               @                       @      @              @      @              �?      @              �?                              @              @                       @                      @              @      M@     �b@      @      K@     �b@               @      @                      �?               @      @               @      @              @      @              �?      �?              �?                              �?              @       @               @       @                      �?               @      �?               @                              �?              @                       @                              �?      @      G@      b@      @      D@     �a@      @      D@     @_@      @      D@     �]@      @      @@      O@      @      1@      3@       @      &@      0@       @      "@      0@       @      @      @       @      �?      @                       @       @      �?      �?              �?               @              �?       @                                      �?              @                      @      *@               @       @                       @               @                       @      &@                       @               @      @                       @               @      �?               @                              �?               @              �?      @      @              �?      @                      @              �?              �?      @              �?       @              �?                               @                      @              @      .@     �E@      @      .@     �@@              ,@      <@                       @              ,@      4@               @      0@              @      ,@               @      @                      @               @                      @      "@                       @              @      �?                      �?              @                       @       @                       @               @                      @      @                      @              @      �?              @      �?              �?      �?              �?                              �?              @                      �?              @      �?      @              �?      @                       @              �?      �?              �?                              �?      @               @      @                                       @                      $@               @      L@              @      &@                      "@              @       @              �?       @              �?                               @              @                      @     �F@                      0@              @      =@              @      "@              �?      �?                      �?              �?                       @       @                      @               @       @              �?       @                       @              �?                      �?                              4@                      @                      0@              @      @                       @              @      �?              @                      @      �?                      �?              @                      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B`         �                    �?T���?�           ��@       �                   �b@�����)�?�            �w@       �                   n@��C,���?�            �s@       ;                   �_@
��F��?�            �j@       .                    �?c�� ��?2            �S@       -                   `_@L)�ڙ�?%            �K@                           W@ZhZ�-�?$            �J@       	                    W@      �?              @������������������������       �                     �?
                          @E@؇���X�?             @                          �\@r�q��?             @������������������������       �                     @                          �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?       (                    �?���Q��?            �F@                          �e@J�fj�?            �B@                          �c@���Q��?             @������������������������       �                     @������������������������       �                      @                           �?      �?             @@                           k@      �?              @                           Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?       !                   `i@r�q��?             8@                           �f@$�q-�?	             *@                          @`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@"       %                     �?���!pc�?             &@#       $                   @\@���Q��?             @������������������������       �                      @������������������������       �                     @&       '                   �a@r�q��?             @������������������������       �                     @������������������������       �                     �?)       *                   �l@      �?              @������������������������       �                     @+       ,                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @/       6                    �?�8��8��?             8@0       3                     �?X�<ݚ�?
             2@1       2                   �Z@���Q��?             @������������������������       �                      @������������������������       �                     @4       5                   �^@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?7       8                   �W@      �?             @������������������������       �                      @9       :                   @_@      �?             @������������������������       �                     @������������������������       �                     �?<       E                    �?\� �D��?S            �`@=       >                     �?<�
I��?             3@������������������������       �                     �??       @                   �b@B{	�%��?
             2@������������������������       �                     (@A       D                    �?VUUUUU�?             @B       C                   `@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @F       g                   @b@�b-�I��?H            �\@G       L                   �`@�G�z�?&             N@H       I                   �_@      �?
             0@������������������������       �                     ,@J       K                   `a@      �?              @������������������������       �                     �?������������������������       �                     �?M       \                    �?fP*L��?             F@N       S                    a@�����?             3@O       R                   `]@���Q��?             @P       Q                   @V@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @T       Y                    �?d}h���?             ,@U       V                    P@�����H�?             "@������������������������       �                     @W       X                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @Z       [                   `]@���Q��?             @������������������������       �                     @������������������������       �                      @]       f                    �?`2U0*��?             9@^       e                   �K@�8��8��?	             (@_       `                     �?ףp=
�?             $@������������������������       �                      @a       d                   �a@      �?              @b       c                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     *@h       }                   �j@|��r��?"             K@i       j                     �?t���]��?             :@������������������������       �                     @k       z                    �?\1�K36�?             7@l       y                   �j@�z�G��?             4@m       r                   �`@      �?
             0@n       q                   �^@�<ݚ�?             "@o       p                   �Z@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @s       x                    �?և���X�?             @t       w                    b@      �?             @u       v                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @{       |                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @~       �                    �?
^N��)�?             <@       �                   `X@�t����?             1@������������������������       �                      @������������������������       �        
             .@�       �                   0l@��!pc�?             &@�       �                   �k@؇���X�?             @������������������������       �                      @�       �                   �^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �l@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �R@&Hk����?D            �Y@������������������������       �                      @�       �                    `@Tt$����?C             Y@�       �                   �X@      �?             @@������������������������       �                     �?�       �                   `p@�g�y��?             ?@�       �                   �`@�C��2(�?             &@������������������������       �                     @�       �                     �?r�q��?             @������������������������       �                     �?�       �                   Hp@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     4@�       �                   Pn@�W��H��?/             Q@������������������������       �                      @�       �                    �?\|/��j�?.            �P@�       �                    d@�n���?             "@�       �                    �?�$I�$I�?             @�       �                   pb@z�G�z�?             @������������������������       �                     @�       �                   q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �p@�MWl��?&            �L@�       �                   pb@�����?             5@������������������������       �                     "@�       �                   `c@r�q��?             (@�       �                   p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@�       �                    �?tk~X��?             B@�       �                   �\@     ��?             @@�       �                   �c@�q�q�?             "@�       �                   q@؇���X�?             @������������������������       �                     @�       �                   @r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   Pa@�㙢�c�?             7@�       �                    b@�IєX�?             1@������������������������       �                     &@�       �                   �w@r�q��?             @�       �                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �a@      �?             @������������������������       �                      @�       �                   �r@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?     0�?'             P@�       �                    p@r-�T��?              J@�       �                   �d@؇���X�?             5@�       �                   �U@@4և���?
             ,@������������������������       �                     �?������������������������       �        	             *@�       �                   �d@����X�?             @������������������������       �                      @������������������������       �                     @�       �                   @c@�Ğ�x��?             ?@�       �                    �?:/����?             <@�       �                     �?��\���?	             1@�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   8r@�θ�?             *@������������������������       �                     @�       �                   Pe@      �?              @�       �                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   `]@"pc�
�?             &@������������������������       �                     @�       �                     �?����X�?             @������������������������       �                     �?�       �                   �q@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �d@��8��8�?             (@�       �                    ^@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       "                   �?���H��?�            @v@�                         �`@@�[�v�?/            @U@�       �                   �^@lJ��?            �H@�       �                   �d@և���X�?             5@�       �                   `V@      �?             0@������������������������       �                     @�       �                   �`@$�q-�?             *@�       �                     �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     @�       �                    �?�m۶m��?             <@�       �                   �e@r�q��?	             2@������������������������       �                     &@�       �                   Pl@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �i@��Q��?             $@������������������������       �                      @�                         Pl@      �?              @                           �?z�G�z�?             @������������������������       �                     �?                         @      �?             @                        ``@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?      
                   �?�q�q�?             @      	                  `o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                        0d@�"e����?             B@                         �?~h����?             <@                        �a@6|���t�?             :@������������������������       �                     &@                        �a@�h$��W�?             .@������������������������       �                     @                          �?�q�q�?             (@������������������������       �                      @                         �?z�G�z�?             $@������������������������       �                     �?                         @�����H�?             "@������������������������       �                     @                        �q@      �?             @                        a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @      !                   @      �?              @                         pi@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @#      J                    �?��Q���?�            �p@$      )                  �\@�yg�;�?4            @R@%      (                   �?      �?             @&      '                  �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?*      I                  q@�㙢�c�?1            @Q@+      :                   �?�θ�?$             J@,      -                  �\@"pc�
�?            �@@������������������������       �                     @.      9                   �?d}h���?             <@/      2                  �^@��+7��?             7@0      1                  �p@�q�q�?             "@������������������������       �                     @������������������������       �                     @3      4                  0`@d}h���?	             ,@������������������������       �                     �?5      6                  �`@8�Z$���?             *@������������������������       �                     @7      8                  �a@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @;      H                   b@�����?             3@<      E                   @��
ц��?
             *@=      B                   �?X�<ݚ�?             "@>      A                  pl@      �?             @?      @                  @_@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @C      D                  �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?F      G                   �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     1@K      t                  �`@(?���?z            �h@L      Y                   �?�����?              O@M      N                  `X@�\��N��?             3@������������������������       �                     @O      T                  �`@     ��?
             0@P      Q                  @_@ףp=
�?             $@������������������������       �                     @R      S                   �?؇���X�?             @������������������������       �                     @������������������������       �                     �?U      X                  `m@      �?             @V      W                  �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @Z      g                   �?L����?            �E@[      `                  �`@$:9$A��?             =@\      ]                  @^@�q�q�?             (@������������������������       �                     @^      _                  �Q@����X�?             @������������������������       �                     @������������������������       �                      @a      f                  c@@�0�!��?             1@b      c                   b@���!pc�?             &@������������������������       �                     @d      e                   _@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @h      o                  `a@~h����?             ,@i      n                   �?؇���X�?             @j      k                  �\@      �?             @������������������������       �                      @l      m                  @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @p      s                   @؇���X�?             @q      r                  �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @u      �                   ]@�H�9��?Z             a@v      {                   �?9��8���?             8@w      x                  �k@      �?              @������������������������       �                     @y      z                  @[@      �?             @������������������������       �                      @������������������������       �                      @|      �                   �?     ��?	             0@}      �                  p@���Q��?             .@~                        Pc@      �?              @������������������������       �                     @�      �                   L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                  `Q@��)x9��?M             \@�      �                   �?�q�q�?             @�      �                   d@���Q��?             @�      �                   `@�q�q�?             @������������������������       �                     �?�      �                  pb@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                   �?�	���?H            �Z@�      �                   �?�Y���U�?>            �V@�      �                  �b@T:�g *�?7            �S@�      �                  pa@     ��?             0@�      �                  �a@d}h���?             ,@������������������������       �                      @�      �                   �?      �?             @�      �                  �a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �                  @g@�=Dފ�?)            �O@�      �                  �m@�ؓo�?(             O@������������������������       �                     ?@�      �                  0e@-���?             ?@�      �                  e@B{	�%��?             2@�      �                  �^@      �?             0@�      �                   d@���Q��?             @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                      @������������������������       �                     *@������������������������       �                     �?�      �                  �p@���|���?             &@�      �                  �c@�<ݚ�?             "@�      �                  o@      �?              @�      �                  pl@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @�      �                   j@      �?
             0@������������������������       �                     *@�      �                  @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KM�KK��h[�B()        K@     �v@     �s@      >@     `o@     @X@      <@     `l@     �M@      *@     �b@     �I@       @      G@      9@      @      ?@      2@      @      ?@      2@      �?      �?      @      �?                              �?      @              �?      @                      @              �?       @              �?                               @                      �?      @      >@      (@      @      =@      @       @      @                      @               @                      �?      :@      @      �?      @      �?              @      �?                      �?              @              �?                              4@      @              (@      �?               @      �?               @                              �?              $@                       @      @              @       @                       @              @                      @      �?              @                              �?              �?      @                      @              �?       @              �?                               @       @                       @      .@      @       @      (@      @       @              @       @                                      @              (@      �?              (@                              �?              @      @                       @              @      �?              @                              �?      @     �Y@      :@       @      .@       @              �?               @      ,@       @              (@               @       @       @       @               @       @                                       @               @              @     �U@      8@      �?      J@      @      �?      .@                      ,@              �?      �?              �?                              �?                     �B@      @              *@      @               @      @               @      �?                      �?               @                               @              &@      @               @      �?              @                       @      �?                      �?               @                      @       @              @                               @              8@      �?              &@      �?              "@      �?               @                      @      �?               @      �?                      �?               @                      @                       @                      *@               @     �A@      1@      �?      &@      ,@              @              �?       @      ,@              @      ,@              @      $@               @      @               @       @                       @               @                              @              @      @              �?      @              �?      �?                      �?              �?                               @              @                              @      �?       @              �?                               @              �?      8@      @              .@       @                       @              .@              �?      "@      �?      �?      @                       @              �?      @              �?                              @                      @      �?                      �?              @              .@     �S@       @       @                      *@     �S@       @              >@       @                      �?              >@      �?              $@      �?              @                      @      �?              �?                      @      �?              @                              �?              4@              *@     �H@      @       @                      &@     �H@      @      @      @       @      �?      @       @              @      �?              @                      �?      �?                      �?              �?              �?              �?      �?                                      �?       @                       @     �F@      @       @      3@                      "@               @      $@               @      �?                      �?               @                              "@              @      :@      @      @      6@      @      @      @              @      �?              @                       @      �?                      �?               @                               @                      3@      @              0@      �?              &@                      @      �?               @      �?               @                              �?              @                      @      @                       @              @      �?                      �?              @                      @               @      8@      C@      �?      2@     �@@              @      2@              �?      *@              �?                              *@               @      @               @                              @      �?      .@      .@      �?      .@      (@      �?      @      $@      �?      @                      @              �?                              @      $@                      @              @      @              @       @                       @              @                              @              "@       @              @                      @       @                      �?              @      �?              @                              �?                      @      �?      @      @              @      @                      @              @              �?               @      �?                                       @      8@     @\@     `k@      @      D@     �C@      @      2@      <@              (@      "@              (@      @                      @              (@      �?              @      �?                      �?              @                      "@                              @      @      @      3@              @      .@                      &@              @      @                      @              @              @      @      @       @                      �?      @      @              �?      @                      �?              �?      @              �?       @              �?                               @                      �?      �?       @              �?      �?                      �?              �?                              �?              @      6@      &@      @      5@      @      @      3@      @              &@              @       @      @      @                               @      @                       @               @       @                      �?               @      �?              @                      @      �?              �?      �?              �?                              �?               @                       @                      �?      @              �?      @              �?                              @                      @      2@     @R@     �f@      �?      ,@      M@      �?       @      �?      �?       @                       @              �?                                      �?              (@     �L@              (@      D@              @      ;@                      @              @      6@              @      1@              @      @                      @              @                      @      &@              �?                       @      &@                      @               @      @                      @               @                              @              @      *@              @      @              @      @              @      @              �?      @              �?                              @               @                      �?       @                       @              �?                       @       @               @                               @                      @                      1@      1@     �M@     �^@      (@      A@      0@      �?      @      (@              @              �?      @      (@      �?              "@                      @      �?              @                      @      �?                              @      @              �?      @                      @              �?                       @              &@      <@      @      @      5@      @      @      @                      @              @       @              @                               @                      ,@      @               @      @              @                      @      @                      @              @                      @              @      @      �?              @      �?              @      �?               @                      �?      �?                      �?              �?                      @              @      �?              @      �?              @                              �?              @                      @      9@     �Z@       @      "@      *@       @              @                      @       @               @                       @       @                              "@      @              "@      @               @      @                      @               @      �?               @                              �?              @                              �?      @      0@     @W@              @       @              @       @              �?       @                      �?              �?      �?              �?                              �?               @                      �?              @      (@     �V@      @      &@      S@      @      @     @Q@              @      &@              @      &@                       @              @      @              �?      @              �?                              @               @                       @              @       @      M@       @       @      M@                      ?@       @       @      ;@       @       @      ,@               @      ,@               @      @               @      �?               @                              �?                       @                      &@       @                                      *@      �?                              @      @               @      @              �?      @              �?       @                       @              �?                              @              �?                       @                      �?      .@                      *@              �?       @                       @              �?        �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�BY         �                   �`@=�C����?�           ��@                          @P@Ff�![��?�            pt@������������������������       �                     @       �                   �s@X8�t-��?�            @t@       d                    �?<N����?�            @r@       a                   P`@�ұ(�b�?{            �h@                           ]@8=���?w             h@                           �?�ങa�?             ?@	                           [@*x9/��?             <@
                           �?VUUUUU�?             "@������������������������       �                     @                          b@      �?             @                          �W@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                           �?ԍx�V�?             3@������������������������       �                     "@                           [@H�z�G�?             $@                          `[@      �?             @������������������������       �                     �?                          `Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           \@      �?             @                          �]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �      �?              @������������������������       �                     @       ^                    s@�]����?a            @d@        '                     �?R7�I���?^            �c@!       $                    �?0�����?             ,@"       #                    `@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@%       &                   @[@�q�q�?             @������������������������       �                      @������������������������       �                     �?(       U                   �p@p�x��?V             b@)       B                    �?�>�5���?L            �_@*       A                   0k@H�w��?1            �U@+       4                    �?������?            �K@,       3                   �j@��-�=��?            �C@-       2                    �?�˹�m��?             C@.       1                    V@�z�G��?             $@/       0                   @_@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     <@������������������������       �                     �?5       @                    d@     ��?	             0@6       ?                   �g@*D>��?             *@7       >                   @b@�g���e�?             &@8       9                    `@B{	�%��?             "@������������������������       �                     �?:       =                    a@      �?              @;       <                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     ?@C       T                    �?~��M��?            �D@D       I                   @c@�������?             8@E       H                   �_@�r����?
             .@F       G                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@J       K                    �?�n���?             "@������������������������       �                     �?L       O                   @Z@      �?              @M       N                   �[@      �?             @������������������������       �                      @������������������������       �                      @P       Q                    [@      �?             @������������������������       �                     �?R       S                   �m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     1@V       Y                   �Z@      �?
             2@W       X                   q@���Q��?             @������������������������       �                     @������������������������       �                      @Z       [                   Hq@�θ�?             *@������������������������       �                      @\       ]                   d@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?_       `                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @b       c                     �?���Q��?             @������������������������       �                      @������������������������       �                     @e       �                    �?�ӽZQ�?9            �W@f       �                   �p@�ء�R�?+            �P@g       v                     �?     @�?!             H@h       u                    �?     @�?	             0@i       p                   �a@�h$��W�?             .@j       o                    `@�<ݚ�?             "@k       n                    ^@�q�q�?             @l       m                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @q       r                    @�q�q�?             @������������������������       �                     @s       t                   `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?w       x                    �?     ��?             @@������������������������       �                     @y       �                   a@N��)x9�?             <@z       {                   �Y@      �?
             0@������������������������       �                     �?|       }                   @^@��S�ۿ?	             .@������������������������       �                     "@~                           _@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             (@�       �                   �b@z�G�z�?             @������������������������       �                      @�       �                   pn@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �j@և���X�?             @�       �                   �U@���Q��?             @������������������������       �                     �?�       �                   @]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?�S����?
             3@�       �                    ]@�θ�?             *@������������������������       �                     @������������������������       �                     $@������������������������       �                     @�       �                   �a@�ٴ��?             ;@�       �                    �?�z�G��?
             4@�       �                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�r����?             .@������������������������       �                      @�       �                   a@����X�?             @������������������������       �                     @������������������������       �                      @�       �                   �e@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @@�       j                  �d@!��+v�?           py@�       �                   �^@     @�?�             s@�       �                   �`@Y�����?            �@@������������������������       �                     @�       �                   `c@���NI�?             =@�       �                    @"pc�
�?             6@�       �                    [@^Cy�5�?             3@�       �                   �a@���I��?             1@�       �                   `b@�q�q�?             @�       �                   a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                   b@      �?              @������������������������       �                     @�       �                    c@�Q����?             @�       �                    �?      �?             @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       I                  �a@%x��K��?�            �p@�       �                   @[@��[~d�?�             l@�       �                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                   �[@2�ҥj��?�            �j@�       �                    �?
;&����?             7@�       �                     �?���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?X�<ݚ�?             2@�       �                   �i@և���X�?
             ,@������������������������       �                     @�       �                   @m@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                   �m@      �?             @������������������������       �                     �?�       �                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     �?�                           �?�q�q��?y             h@�                         �`@���,(�?P            �_@�       �                    a@j#�t�?5            �T@������������������������       �                      @�                         ``@���A*��?4            @T@�       �                   i@�MLq��?.            �P@�       �                   Pf@;�;��?	             *@�       �                   e@���Q��?             @������������������������       �                      @�       �                   �e@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �h@      �?              @�       �                    �?�q�q�?             @�       �                     �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   hp@�{��?��?%             K@�       �                   �m@؇���X�?             <@�       �                     �?�<ݚ�?             2@������������������������       �                      @�       �                   0m@���Q��?             $@�       �                    �?      �?              @������������������������       �                      @�       �                    l@�q�q�?             @�       �                   �^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     $@�                          d@R�}e�.�?             :@�                           �?��Q��?             4@�       �                    ]@z�G�z�?             $@������������������������       �                      @�       �                    �?      �?              @�       �                    `@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   0u@�q�q�?             @������������������������       �                     �?������������������������       �                      @      
                   �?      �?             $@      	                  �b@X�<ݚ�?             "@                         �?r�q��?             @                        @_@      �?             @������������������������       �                      @                        `a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@                          �?�eP*L��?             F@                        �a@����X�?             ,@������������������������       �                     @                         �?�C��2(�?             &@                        �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                         �?�q�q�?             >@                         �?�θ�?             :@                        @a@���!pc�?             6@������������������������       �                     @                         �?�����H�?             2@������������������������       �                     �?                        �`@�t����?             1@������������������������       �                      @������������������������       �        
             .@������������������������       �                     @������������������������       �                     @!      (                  Pa@�NoS{�?)            @P@"      '                   �?ףp=
�?             4@#      $                    �?�}�+r��?             3@������������������������       �                     @%      &                  q@��S�ۿ?
             .@������������������������       �        	             ,@������������������������       �                     �?������������������������       �                     �?)      4                  pb@�L�lRT�?            �F@*      /                   �?�t����?
             1@+      .                   �?�q�q�?             @,      -                   b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?0      1                  �o@@4և���?             ,@������������������������       �                     (@2      3                  �`@      �?              @������������������������       �                     �?������������������������       �                     �?5      D                   d@:/����?             <@6      C                   `@;n,�R�?             6@7      <                   �?���Q��?             .@8      9                   ^@      �?             @������������������������       �                      @:      ;                  �_@      �?              @������������������������       �                     �?������������������������       �                     �?=      @                  p@���|���?             &@>      ?                  Ph@r�q��?             @������������������������       �                     �?������������������������       �                     @A      B                  �]@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @E      H                  @l@r�q��?             @F      G                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @J      _                   �?Z��D�?             G@K      ^                   �?ӧ
�.�?             ?@L      S                  �b@Y��sd�?             =@M      R                  �c@����X�?             ,@N      O                  0b@r�q��?             (@������������������������       �                     "@P      Q                  8p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @T      Y                   �?�q�q�?
             .@U      V                   c@      �?              @������������������������       �                     @W      X                  �q@z�G�z�?             @������������������������       �                     �?������������������������       �                     @Z      [                  `c@؇���X�?             @������������������������       �                     @\      ]                  @n@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @`      g                  `c@N贁N�?             .@a      b                  �b@z�G�z�?             $@������������������������       �                     @c      f                   �?����X�?             @d      e                   g@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?h      i                  pd@���Q��?             @������������������������       �                      @������������������������       �                     @k      �                   �?">�Tr^�?E            �Y@l      y                    �?\�r�<,�?>            �V@m      n                  �b@8�Z$���?             :@������������������������       �                      @o      p                  �i@�8��8��?             8@������������������������       �                     &@q      x                  �`@8�Z$���?	             *@r      u                   �?"pc�
�?             &@s      t                  �]@      �?              @������������������������       �                     �?������������������������       �                     �?v      w                  �j@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @z      �                   @nk���L�?-            @P@{      |                  pl@�G�z��?+             N@������������������������       �                     <@}      �                  `]@     ��?             @@~      �                  hp@������?             @      �                  �m@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                   �?HP�s��?             9@�      �                  �^@���N8�?             5@�      �                  0e@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             0@�      �                   q@      �?             @�      �                  �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                  0f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                   �?VUUUUU�?             (@�      �                  �Z@z�G�z�?             @�      �                   f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B(&       �I@     �w@     0s@      @@     �l@      P@                      @      @@     �l@     �N@      @@     �h@     �N@      7@     �b@      9@      7@     �b@      6@      @      2@      @      @      2@      @      @      @      @                      @      @      @              �?      @                      @              �?                       @                      @      .@      �?              "@              @      @      �?              @      �?              �?                       @      �?                      �?               @              @      @               @       @               @                               @              �?      �?                              @      1@     @`@      .@      .@      `@      .@       @      $@       @              $@      �?                      �?              $@               @              �?       @                                      �?      *@     �]@      *@      $@     �Z@      $@       @     @R@      @       @      E@      @      @     �A@              @     �A@              @      @              @       @              @                               @                      @                      <@              �?                      @      @      @      �?      @      @      �?      @      @      �?      @      �?      �?                              @      �?              �?      �?              �?                              �?              @                               @                       @      @                              ?@               @      A@      @       @      1@      @              *@       @              �?       @              �?                               @              (@               @      @      @                      �?       @      @       @               @       @               @                               @       @       @                      �?               @      �?               @                              �?                      1@              @      (@      @      @       @              @                               @                      $@      @                       @              $@      �?              $@                              �?       @      �?                      �?               @                               @      @               @                              @      "@     �H@      B@      @     �@@      ?@      @      >@      .@       @      @      @       @      @      @              @       @              �?       @              �?      �?              �?                              �?                      �?              @               @              @                      @       @              �?       @                                      �?                      �?      �?      7@       @              @              �?      3@       @      �?      ,@      �?                      �?      �?      ,@                      "@              �?      @              �?                              @                      @      @              �?      @                       @              �?       @                       @              �?                      @      @               @      @              �?                      �?      @                      @              �?                       @                      @      0@              @      $@              @                              $@                      @      @      0@      @      @      ,@              @      �?              @                              �?               @      *@                       @               @      @                      @               @                               @      @                      @               @                      @@              3@      b@     `n@      .@     �_@     @d@      @      3@      $@                      @      @      3@      @      @      (@      @      @      "@      @      @      @      @              @       @              �?       @              �?                               @              @              @      @      @      @                      �?      @      @                      @      �?      @      �?      �?      @              �?       @              �?                               @                      �?                              �?               @                      @                      @              &@      [@      c@      @     �T@     @a@              �?      "@              �?                              "@      @     @T@      `@              (@      &@               @      @                       @               @      �?              �?      �?              �?                              �?              �?                      $@       @               @      @              @                      @      @                      @              @                       @       @              �?                      �?       @                       @              �?              @     @Q@     �]@      @     �B@     �U@      @      1@      O@       @                       @      1@      O@       @      1@      H@       @      @      @       @              @                       @       @              �?       @                                      �?              @       @              @       @              �?       @              �?                               @              @                       @                      &@     �E@              @      8@              @      ,@                       @              @      @               @      @                       @               @      @               @       @                       @               @                               @               @                              $@              @      3@              @      *@               @       @                       @               @      @              �?      @                      @              �?                      �?       @              �?                               @              @      @              @      @              �?      @              �?      @                       @              �?      �?              �?                              �?                       @              @                      �?                              @                      ,@              4@      8@              $@      @                      @              $@      �?               @      �?               @                              �?               @                      $@      4@              @      4@              @      0@              @                       @      0@                      �?               @      .@               @                              .@                      @              @              �?      @@      @@               @      2@              �?      2@                      @              �?      ,@                      ,@              �?                      �?              �?      >@      ,@              .@       @               @      �?              �?      �?                      �?              �?                      �?                      *@      �?              (@                      �?      �?                      �?              �?              �?      .@      (@      �?      $@      &@      �?      $@      @      �?      @                       @              �?      �?              �?                              �?                      @      @              @      �?                      �?              @                       @      @                      @               @                              @              @      �?               @      �?                      �?               @                      @              @      :@      ,@      @      .@      (@      @      .@      $@      @      $@               @      $@                      "@               @      �?               @                              �?               @                              @      $@              @      @              @                      �?      @              �?                              @              �?      @                      @              �?      @                      @              �?                               @       @      &@       @       @       @                      @               @      @               @      @                      @               @                              �?                      @       @                       @              @              @      2@     @T@      @      &@     @S@              @      6@               @                       @      6@                      &@               @      &@               @      "@              �?      �?                      �?              �?                      �?       @              �?                               @                       @      @      @     �K@      @      @      K@                      <@      @      @      :@      �?      @      @      �?              @      �?                                      @              @               @              7@      �?              4@      �?              @      �?                                      @                      0@      �?              @      �?              �?      �?                                      �?                       @              @      �?              @                              �?      �?      @      @      �?              @      �?              �?                      �?      �?                                      @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B8i         b                     �?��K��?�           ��@       W                    �?hQ��?]            @a@                          �Z@���Ȅ�?Q            �]@������������������������       �                     @                           �?����2b�?L            @\@                           `@t�����?            �A@                          `T@@�0�!��?
             1@������������������������       �                     �?	       
                   �\@      �?	             0@������������������������       �                     @                           �?�<ݚ�?             "@������������������������       �                     @                           �?�q�q�?             @                          �p@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?B{	�%��?             2@                          �c@h/�����?             "@                          c@r�q��?             @������������������������       �                     @������������������������       �                     �?                          d@�q�q�?             @                          `o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@       "                   �\@��\���?5            �S@        !                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?#       .                    �?�+e�X�?3            �R@$       %                   �b@���Q��?             .@������������������������       �                     @&       -                   �`@�eP*L��?             &@'       (                   `o@����X�?             @������������������������       �                     �?)       ,                   pd@r�q��?             @*       +                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @/       <                    �?z�G�z�?(             N@0       5                   �^@�t����?             A@1       2                   �p@z�G�z�?             $@������������������������       �                     @3       4                    q@�q�q�?             @������������������������       �                      @������������������������       �                     �?6       7                   �`@�8��8��?             8@������������������������       �                     ,@8       ;                   �q@z�G�z�?             $@9       :                   �i@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @=       >                   @Z@�	j*D�?             :@������������������������       �                     @?       J                   �j@���|���?             6@@       I                    @X�<ݚ�?             "@A       B                   �Q@      �?              @������������������������       �                     �?C       H                   �_@����X�?             @D       E                   �\@r�q��?             @������������������������       �                     �?F       G                    b@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?K       V                    @�θ�?	             *@L       S                   �_@      �?             (@M       R                   �^@�����H�?             "@N       O                    k@      �?              @������������������������       �                     @P       Q                   �n@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?T       U                   c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?X       ]                   �^@$����%�?             3@Y       Z                   �Z@���Q��?             @������������������������       �                      @[       \                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?^       _                   �`@����X�?	             ,@������������������������       �                     @`       a                   �p@���Q��?             $@������������������������       �                     @������������������������       �                     @c       �                   �?8l�����?y           ��@d       3                  �b@������?'           p}@e       �                   �`@P�]��k�?�            �s@f       i                   �Q@�a!�z��?}            �h@g       h                   �`@      �?             @������������������������       �                      @������������������������       �                      @j       q                   �X@z���ڜ�?{            @h@k       p                   �U@(;L]n�?             >@l       m                    V@�8��8��?             (@������������������������       �                      @n       o                    b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@r       �                    �?$�*���?j            �d@s       ~                    [@�ȭ����?K            @^@t       u                    �?��\���?             1@������������������������       �                      @v       w                   �\@���Q��?	             .@������������������������       �                     @x       }                    �?�C��2(�?             &@y       |                    X@؇���X�?             @z       {                   �Z@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       �                   @^@�g\��?@             Z@�       �                   �_@�L���?            �B@�       �                   �\@Pa�	�?            �@@�       �                    �?��S�ۿ?             .@������������������������       �                     @�       �                   p`@      �?              @�       �                   `\@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �        
             2@�       �                    `@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?���Ƨ��?-            �P@�       �                   b@r�qG�?             H@�       �                   �]@��� =�?             A@�       �                   0a@      �?
             0@������������������������       �                     "@�       �                   �a@؇���X�?             @�       �                   �g@r�q��?             @������������������������       �                     @�       �                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �^@r�q��?             2@������������������������       �                     �?�       �                   �_@�t����?             1@�       �                   @j@�<ݚ�?             "@�       �                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   pb@�$I�$I�?	             ,@������������������������       �                      @�       �                   �[@�q�q�?             (@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?E�ϣ1��?             3@������������������������       �                     @�       �                   �_@ƒ_,���?             .@������������������������       �                     @�       �                   @c@      �?
             (@�       �                   @a@����X�?             @������������������������       �                     @�       �                    ^@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �d@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    a@���{�?            �E@�       �                   @L@��WV��?	             *@�       �                    _@��8��8�?             (@�       �                    _@B{	�%��?             "@������������������������       �                     �?�       �                    �?      �?              @������������������������       �                      @�       �                    �?r�q��?             @�       �                   @]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    `@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?d��0u��?             >@�       �                   @_@"pc�
�?             &@�       �                   �Z@���Q��?             @�       �                   �k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   `^@�\��N��?             3@�       �                    @���!pc�?             &@�       �                   �j@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   `]@      �?              @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �[@p=
ףp�?M             ^@�       �                    �?     ��?
             0@������������������������       �                     (@�       �                    �?      �?             @�       �                   m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       "                  �a@8�Z$���?C             Z@�                         �a@TQm�y�?3            �R@�       �                    �?�[�IJ�?            �G@�       �                   �p@��S�r
�?             <@�       �                   �_@�G�z�?             4@�       �                   �^@      �?              @�       �                   �h@�q�q�?             @������������������������       �                     @�       �                    o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   �j@      �?             (@�       �                    �?      �?             @�       �                    �?���Q��?             @�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   @_@      �?              @������������������������       �                     @�       �                   8s@���Q��?             @������������������������       �                     @������������������������       �                      @�                          �?�KM�]�?             3@�                         r@�r����?
             .@�                          0i@@4և���?	             ,@�       �                   Pa@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?������������������������       �                     @                         �?Dc}h��?             <@������������������������       �                      @      !                   @t���]��?             :@                         0a@�^)��?             9@                        �g@;n,�R�?             6@	                         T@p=
ףp�?             $@
                        @_@      �?              @������������������������       �                     �?������������������������       �                     �?                         �?      �?              @                        �b@      �?             @                        @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @                        �j@      �?
             (@������������������������       �                     @                         l@�q�q�?             "@������������������������       �                     �?                         b@      �?              @������������������������       �                      @                        �b@�q�q�?             @������������������������       �                     �?                         �?z�G�z�?             @������������������������       �                      @                        0m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?#      2                   �?^ev��?             =@$      /                  0q@     @�?             0@%      .                   �?p=
ףp�?             $@&      -                   �?B{	�%��?             "@'      (                   �?      �?             @������������������������       �                     @)      *                  �b@VUUUUU�?             @������������������������       �                     �?+      ,                  �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?0      1                  �s@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     *@4      y                   @@��-�=�?]             c@5      d                  �p@>N&� �?X             b@6      S                   �?�X���?A             \@7      @                  i@��ż1�?,            @S@8      ?                  �d@�GN�z�?             6@9      >                  �h@�eP*L��?             &@:      ;                  Pd@      �?              @������������������������       �                     @<      =                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@A      B                  �k@����n��?             �K@������������������������       �                     6@C      D                  d@��!pc�?            �@@������������������������       �                     &@E      H                  �\@�X����?             6@F      G                   f@���Q��?             @������������������������       �                     @������������������������       �                      @I      R                   �?@�0�!��?             1@J      Q                  �n@      �?
             0@K      N                   �?���Q��?             @L      M                  0a@�q�q�?             @������������������������       �                     �?������������������������       �                      @O      P                  `f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?T      Y                  pc@��Ħ��?            �A@U      X                  0n@��!pc�?             &@V      W                   �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @Z      a                   �?r�q��?             8@[      `                   �?�KM�]�?             3@\      ]                  `l@�q�q�?             @������������������������       �                     �?^      _                   `@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     *@b      c                  @e@���Q��?             @������������������������       �                     @������������������������       �                      @e      f                  0c@���|���?            �@@������������������������       �                     @g      n                   �?X�<ݚ�?             ;@h      m                  �r@�q�q�?             (@i      j                  @_@      �?              @������������������������       �                     @k      l                  �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @o      t                   �?�q�q�?             .@p      s                  @`@����X�?             @q      r                  s@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @u      x                  u@      �?              @v      w                  �p@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @z      {                  d@      �?              @������������������������       �                     @|      }                   �?�q�q�?             @������������������������       �                     �?~                         �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  P`@�z�΅�?R            @_@�      �                  �j@+�W�?8            �U@�      �                   `@�2(&��?             F@�      �                  j@��WV��?            �C@�      �                   �?�3�2%��?            �A@�      �                   �?r�q��?             8@�      �                   �?��#��Z�?             6@�      �                  @U@��8��8�?
             (@�      �                  �^@���(\��?             $@������������������������       �                      @�      �                  `]@      �?              @������������������������       �                     @�      �                  @^@�Q����?             @�      �                  �]@      �?             @������������������������       �                     �?�      �                  P`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �                  `^@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                      @�      �                   �?�eP*L��?             &@������������������������       �                     @�      �                   @����X�?             @�      �                  �]@�q�q�?             @������������������������       �                      @�      �                   ^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   �?�Q����?             @�      �                  �b@      �?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                  @^@AA�?             E@�      �                   ]@���Q��?             @�      �                   Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �                  �o@@0.1�r�?            �B@������������������������       �                     4@�      �                   `@�"�O�|�?             1@�      �                   �?��S�ۿ?             .@�      �                  �]@ףp=
�?             $@������������������������       �                     @�      �                  �e@      �?             @������������������������       �                     �?�      �                  �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�      �                  ``@�99lMt�?            �C@�      �                  pe@      �?             0@�      �                   �?����X�?             ,@�      �                   �?؇���X�?             @�      �                  �m@      �?             @������������������������       �                      @�      �                  �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                  Pb@և���X�?             @�      �                  �g@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �_@      �?             @�      �                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                  @a@�㙢�c�?             7@������������������������       �                     @�      �                  �a@������?
             1@�      �                  pb@���Q��?             @�      �                  �a@      �?             @�      �                   Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�      �                   a@�8��8��?             (@������������������������       �                     @�      �                   �?z�G�z�?             @�      �                  b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B-       �I@     �v@     t@      @     �J@     �S@      @     �E@     @R@              @              @     �B@     @R@       @      1@      0@              @      ,@              �?                       @      ,@                      @               @      @                      @               @      @              �?       @                       @              �?                      �?       @                       @              �?               @      ,@       @       @      @       @      �?      @                      @              �?                      �?               @      �?              �?                      �?      �?                                      �?              "@              �?      4@     �L@      �?       @                       @              �?                              2@     �L@              @      "@                      @              @      @               @      @              �?                      �?      @              �?       @                       @              �?                              @              @                      (@      H@              @      >@               @       @                      @               @      �?               @                              �?               @      6@                      ,@               @       @               @       @                       @               @                              @               @      2@                      @               @      ,@              @      @              @      @                      �?              @       @              @      �?              �?                      @      �?                      �?              @                              �?                      �?              @      $@              @      "@              �?       @              �?      @                      @              �?      @              �?                              @                      �?               @      �?               @                              �?                      �?      @      $@      @      @               @       @                      �?               @                       @      �?                              $@      @              @                      @      @              @                              @     �F@     Ps@     @n@      A@     �m@      i@      ;@      i@     �V@      5@     �a@      B@       @               @       @                                       @      3@     �a@      A@      �?      =@              �?      &@                       @              �?      @                      @              �?                              2@              2@      \@      A@      ,@     �W@      *@      @      $@      �?       @                      @      $@      �?      @                              $@      �?              @      �?              @      �?              @                              �?              @                      @               @      U@      (@      @      A@              �?      @@              �?      ,@                      @              �?      @              �?      @                      @              �?                               @                      2@               @       @               @                               @              @      I@      (@      @      C@      @      �?      >@      @      �?      .@                      "@              �?      @              �?      @                      @              �?       @                       @              �?                              �?                      .@      @                      �?              .@       @              @       @              �?       @              �?                               @              @                       @               @       @      @       @                               @      @               @      @                      @               @                      @               @      (@      @              @               @       @      @                      @       @       @       @              @       @              @                       @       @               @                               @       @      @               @                              @              @      2@      5@      @      @       @      @      @       @      �?      @      �?      �?                              @      �?               @                      @      �?               @      �?                      �?               @                      @               @              �?       @                                      �?      �?                              &@      3@               @      "@               @      @               @      �?                      �?               @                               @                      @              "@      $@               @      @              @      @                      @              @                       @                      �?      @              �?      �?                      �?              �?                              @      @      N@      K@              *@      @              (@                      �?      @              �?      �?                      �?              �?                               @      @     �G@     �I@      @      <@      F@       @      .@      >@       @      *@      *@       @      &@      @       @       @      @               @      @                      @               @      �?               @                              �?       @                              "@      @              @      @              @       @               @       @               @                               @              �?                              �?              @                       @      @                      @               @      @                      @               @                       @      1@               @      *@              �?      *@              �?      @                      @              �?                              $@              �?                              @      �?      *@      ,@               @              �?      &@      ,@      �?      $@      ,@      �?      $@      &@      �?      @       @              �?      �?                      �?              �?              �?      @      �?      �?       @      �?      �?              �?      �?                                      �?               @                      @                      @      "@                      @              @      @              �?                       @      @                       @               @      @              �?                      �?      @                       @              �?       @                       @              �?                              @              �?              @      3@      @      @      @      @      �?       @      @      �?      �?      @      �?      �?      @                      @      �?      �?      �?      �?                              �?      �?                      �?              �?                              @              �?               @      @                      @               @                              *@              @      B@     �[@      @      =@     @[@      @      1@      V@      @       @     �P@              @      1@              @      @               @      @                      @               @      �?               @                              �?              @                              &@      @      @     �H@                      6@      @      @      ;@                      &@      @      @      0@      @               @      @                                       @              @      ,@               @      ,@               @      @              �?       @              �?                               @              �?      �?                      �?              �?                              &@              �?              @      "@      6@      @      @       @      @      @                      @              @                                       @              @      4@               @      1@               @      @                      �?               @      @               @                              @                      *@               @      @                      @               @                      (@      5@                      @              (@      .@              @      @              @      �?              @                      @      �?                      �?              @                              @              @      $@               @      @               @      �?               @                              �?                      @              @      @              �?      @              �?                              @               @                      @      �?              @                       @      �?              �?                      �?      �?                      �?              �?              &@      R@      E@      &@      M@      1@      "@      6@      *@      @      5@      (@      @      5@       @      �?      .@       @      �?      .@      @      �?      @      @      �?      @      @                       @      �?      @      @              @              �?      �?      @      �?              @                      �?      �?               @      �?                                       @              �?                       @                      "@      �?                      �?              "@                               @      @      @                      @              @       @              @       @               @                       @       @               @                               @              �?                                      @      @      �?      �?      @      �?              �?      �?                      �?              �?                       @                                      �?       @      B@      @               @      @               @      �?                      �?               @                               @       @      A@      �?              4@               @      ,@      �?              ,@      �?              "@      �?              @                      @      �?              �?                       @      �?                      �?               @                      @               @                              ,@      9@              $@      @              $@      @              @      �?              @      �?               @                      �?      �?                      �?              �?                      @                      @      @               @      �?                      �?               @                       @       @              �?       @                       @              �?                      �?                               @              @      3@                      @              @      *@              @       @              @      �?               @      �?                      �?               @                      �?                              �?              �?      &@                      @              �?      @              �?      �?              �?                              �?                      @�t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�_         N                  �c@��J��?�           ��@       �                   `@�P����?d           ��@       n                    �?����?�            �q@       ;                    `@"�l0��?�            �i@                           �[@/y0��k�?0            �S@                          �h@     ��?             @@                           �?�n���?
             2@       	                   �Y@�8��8��?             (@������������������������       �                     @
                          `_@�n���?             "@������������������������       �                     @                          �_@���Q��?             @������������������������       �                      @������������������������       �                     @                          �^@VUUUUU�?             @                           �?      �?             @                          @Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @                          �Y@0�����?             ,@������������������������       �                     @                          �Y@h/�����?             "@������������������������       �                      @                           �?����X�?             @������������������������       �                      @                           �?���Q��?             @                          pn@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?!       ,                    �?K����?             G@"       +                   `_@6YE�t�?            �@@#       $                     �?��S�ۿ?             >@������������������������       �                     �?%       *                    �? 	��p�?             =@&       )                   Po@      �?              @'       (                   �^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     5@������������������������       �                     @-       8                    �?;�;��?	             *@.       /                     �?�n���?             "@������������������������       �                     �?0       1                   �Z@      �?              @������������������������       �                     @2       7                    ^@�Q����?             @3       4                   `\@      �?             @������������������������       �                      @5       6                   @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?9       :                    _@      �?             @������������������������       �                     �?������������������������       �                     @<       G                   �O@�8ui�?X            �_@=       B                   `]@b�h�d.�?            �A@>       A                   0a@���N8�?             5@?       @                   �Q@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     (@C       D                    �?X�Cc�?             ,@������������������������       �                     @E       F                   @^@����X�?             @������������������������       �                     @������������������������       �                      @H       a                    �?������?B            �V@I       V                    a@     ��?/             P@J       U                    �?�(\����?             4@K       P                   �`@�"�O�|�?             1@L       M                   pm@@4և���?
             ,@������������������������       �                     $@N       O                   �X@      �?             @������������������������       �                     �?������������������������       �                     @Q       R                   �`@VUUUUU�?             @������������������������       �                     �?S       T                   �o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @W       `                   0k@���7�?              F@X       _                   k@"pc�
�?             &@Y       Z                   pe@ףp=
�?             $@������������������������       �                     @[       ^                    �?z�G�z�?             @\       ]                   Pg@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                    �@@b       m                   �\@�+$�jP�?             ;@c       l                   �[@X�Cc�?
             ,@d       g                    �?"pc�
�?             &@e       f                   `b@      �?              @������������������������       �                     �?������������������������       �                     �?h       k                    a@�����H�?             "@i       j                   �t@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        	             *@o       �                    `@�_�(�?5            �S@p       �                    �?��(\���?             4@q       v                    �?�S����?             3@r       s                   `]@r�q��?             @������������������������       �                     @t       u                    @      �?              @������������������������       �                     �?������������������������       �                     �?w       z                    �?��WV��?
             *@x       y                   �^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @{       �                   �U@      �?              @|       }                   �W@      �?             @������������������������       �                     �?~                          `\@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �[@      �?             @�       �                   r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?*Շ�b�?&            �M@�       �                   �X@t����{�?            �B@������������������������       �                     @�       �                   c@z5�h$�?             >@�       �                   @a@z�G�z�?             @�       �                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   pb@tF��_�?             9@�       �                     �?�d�����?             3@������������������������       �                     @�       �                    �?     ��?
             0@������������������������       �                     @�       �                    �?�eP*L��?             &@�       �                    �?X�<ݚ�?             "@������������������������       �                     @�       �                   `_@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �\@r�q��?             @�       �                   pk@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   `\@8�A�0��?             6@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?	             (@�       �                   �a@�8��8��?             @�       �                    _@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �X@r�q��?             @������������������������       �                     �?������������������������       �                     @�                          �?8s���?�            Pq@�       �                   0g@�+78�/�?S            �a@�       �                   Pa@x��s���?            �D@�       �                    �? )O��?             B@�       �                     �?j���� �?             1@������������������������       �                     @�       �                   �`@�q�q�?             (@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                    a@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   `]@�˹�m�?             3@�       �                     �?      �?              @������������������������       �                     �?�       �                   Pa@����X�?             @�       �                   @Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                    �?z�G�z�?             @�       �                   �e@      �?             @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?�EL�o�?:            �X@�       �                    �?�������?0            @T@�       �                   �s@�
���?)            �P@�       �                   �_@2�����?#             K@�       �                    c@
ףp=
�?             4@�       �                   @b@�˹�m�?             3@�       �                   �p@�.�?��?
             .@�       �                   �j@�؉�؉�?	             *@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �\@��(\���?             $@�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �^@      �?              @������������������������       �                     @�       �                   `k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   Pc@l��\��?             A@�       �                     �?      �?             @@������������������������       �                     (@�       �                   �l@P���Q�?             4@�       �                   c@r�q��?             @������������������������       �                     @�       �                   �f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             ,@������������������������       �                      @�       �                   �t@�q�q�?             (@������������������������       �                     @������������������������       �                     @�       �                     �?���Q��?             .@������������������������       �                     �?�       �                   `c@����S�?             ,@�       �                   `p@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                     �?�                         `a@�)O�?
             2@�       �                     �?      �?             @������������������������       �                     �?�       �                   Pn@VUUUUU�?             @������������������������       �                     �?                         t@      �?              @������������������������       �                     �?������������������������       �                     �?                        �e@؇���X�?             ,@������������������������       �                     (@������������������������       �                      @                         �?�j��z�?T             a@                        pa@�{��?��?"             K@                        0p@�˹�m��?             C@	                         �?�S����?             3@
                        �^@d}h���?             ,@                        p@�����H�?             "@������������������������       �                      @������������������������       �                     �?                        b@���Q��?             @                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �        	             3@                        hp@      �?
             0@������������������������       �                     @                        a@���!pc�?             &@������������������������       �                      @                        �q@�����H�?             "@                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @      M                  0b@�X�=ٚ�?2            �T@      4                  pl@b�*j��?+            @R@       /                   �?��\Wن�?             =@!      "                    �?�GN�z�?             6@������������������������       �                      @#      .                  Pc@      �?             4@$      -                  �`@r�q��?             2@%      *                   �?�t����?             1@&      )                  �g@�8��8��?             (@'      (                   g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@+      ,                  Pa@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @0      1                  �g@:/����?             @������������������������       �                     @2      3                  �i@      �?             @������������������������       �                      @������������������������       �                      @5      L                   �?5_�g���?             F@6      ?                  b@�p\�y�?            �D@7      >                  0a@      �?	             4@8      =                  Xr@�q�q�?             (@9      :                   @�<ݚ�?             "@������������������������       �                     @;      <                  �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @@      A                  �b@ܤ�[r�?             5@������������������������       �                      @B      C                  �b@/y0��k�?	             *@������������������������       �                     @D      K                  p`@      �?              @E      J                  �^@�8��8��?             @F      G                  �Z@�q�q�?             @������������������������       �                     �?H      I                  pm@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     $@O      v                   �?lYVn�?k            �e@P      u                  �f@Rg��J��?            �H@Q      l                  �q@��6���?             E@R      _                    �?     ��?             @@S      ^                   �?�eP*L��?	             &@T      ]                  hp@      �?             $@U      V                  �`@����X�?             @������������������������       �                      @W      \                  Pe@���Q��?             @X      [                  d@      �?             @Y      Z                  �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?`      k                   �?���N8�?             5@a      b                   �?�d�����?             3@������������������������       �                      @c      h                  Pe@@�0�!��?	             1@d      e                  pd@$�q-�?             *@������������������������       �                     @f      g                  �a@      �?              @������������������������       �                     @������������������������       �                     �?i      j                   n@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @m      t                   �?z�G�z�?             $@n      o                  �r@����X�?             @������������������������       �                     �?p      q                  �`@r�q��?             @������������������������       �                     @r      s                  �u@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @w      x                  �c@6_%��?L            @_@������������������������       �                     "@y      �                  �^@��6�8�?I             ]@z      �                  f@,�����?             �H@{      �                   �?���
�?            �A@|      �                  �e@�g���e�?            �@@}      �                  @i@N��)x9�?             <@~                        �X@      �?             @������������������������       �                      @�      �                  �Z@      �?             @������������������������       �                     �?������������������������       �                     @�      �                  �d@�GN��?             6@�      �                   �?�����H�?             "@������������������������       �                     @�      �                  �o@z�G�z�?             @������������������������       �                     @�      �                  �\@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?8�Z$���?	             *@�      �                  e@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �d@p=
ףp�?             $@������������������������       �                      @�      �                   m@      �?              @������������������������       �                     @�      �                  �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                  �r@؇���X�?
             ,@������������������������       �        	             (@������������������������       �                      @�      �                   �?t�U����?)            �P@�      �                  �`@ �h�7W�?             �J@������������������������       �        
             3@�      �                  a@l��\��?             A@�      �                  d@�q�q�?             @������������������������       �                      @�      �                    @      �?             @������������������������       �                      @������������������������       �                      @�      �                   b@h�����?             <@�      �                  �d@�IєX�?	             1@������������������������       �                     �?������������������������       �                     0@������������������������       �        	             &@�      �                  po@X�Cc�?	             ,@�      �                  �d@X�<ݚ�?             "@�      �                    �?և���X�?             @������������������������       �                     �?�      �                   �?�q�q�?             @�      �                  �d@      �?             @������������������������       �                     �?������������������������       �                     @�      �                  �U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B�(        H@     0x@     �r@     �G@     Pu@     �e@     �A@     @h@      K@      :@     �c@      4@      2@      H@      (@       @      ,@      $@      @      @       @      @       @      @                      @      @       @      @      @                               @      @               @                              @       @       @       @       @       @               @      �?                      �?               @                              �?                               @       @      $@       @              @               @      @       @                       @       @      @                       @               @      @               @       @                       @               @                              �?              $@      A@       @      @      <@               @      <@                      �?               @      ;@               @      @               @       @                       @               @                              @                      5@              @                      @      @       @      @      @       @                      �?      @      @      �?      @                      �?      @      �?      �?      @                       @              �?      �?              �?                              �?                              �?      �?      @              �?                              @               @     �[@       @              =@      @              4@      �?               @      �?                      �?               @                      (@                      "@      @              @                       @      @                      @               @               @     @T@       @      @     �M@       @      �?      1@       @      �?      ,@       @              *@      �?              $@                      @      �?                      �?              @              �?      �?      �?      �?                              �?      �?                      �?              �?                      @               @      E@               @      "@              �?      "@                      @              �?      @              �?      �?              �?                              �?                      @              �?                             �@@              @      6@              @      "@               @      "@              �?      �?              �?                              �?              �?       @              �?      �?                      �?              �?                              @              @                              *@              "@      B@      A@      @      @      (@      @      @      (@      �?              @                      @      �?              �?      �?                                      �?       @      @      @              �?      @              �?                              @       @      @      @       @       @                      �?               @      �?                      �?               @                              �?      @              �?      �?                      �?              �?                               @              �?              @      ?@      6@       @      0@      3@              @               @      "@      3@      �?      @              �?      �?                      �?              �?                              @              �?      @      3@              @      ,@                      @              @      &@                      @              @      @              @      @                      @              @       @              @                               @              �?      �?              �?                              �?      �?              @      �?              �?                      �?      �?                                      @      @      .@      @      �?      "@                      @              �?       @              �?                               @              @      @      @       @      �?      @       @      �?               @                              �?                              @      �?      @              �?                              @              (@     `b@     �]@      @     @Y@      @@       @      7@      0@      �?      7@      (@              $@      @              @                      @      @                      @              @      @              @                       @      @               @                              @      �?      *@      @      �?       @      @      �?                               @      @               @      �?               @                              �?                      @              &@              �?              @      �?              @      �?              �?      �?                                      �?                       @                      �?      @     �S@      0@       @      P@      .@      �?     �I@      ,@      �?      F@      "@      �?      *@      @      �?      *@      @      �?      "@      @      �?      "@      @              �?       @                       @              �?              �?       @      �?              �?      �?              �?                              �?      �?      @                      @              �?      �?                      �?              �?                                       @              @                              �?              ?@      @              ?@      �?              (@                      3@      �?              @      �?              @                      �?      �?                      �?              �?                      ,@                               @              @      @                      @              @              �?      *@      �?              �?              �?      (@      �?              (@      �?              (@                              �?      �?                      @      ,@      �?      �?       @      �?              �?              �?      �?      �?                      �?      �?      �?              �?                              �?               @      (@                      (@               @                      @      G@     �U@              &@     �E@              @     �A@              @      0@              @      &@              �?       @                       @              �?                       @      @               @      �?                      �?               @                               @                      @                      3@               @       @                      @               @      @                       @               @      �?              �?      �?                      �?              �?                      @              @     �A@     �E@      @      9@     �E@       @      @      4@              @      1@                       @              @      .@              @      .@               @      .@              �?      &@              �?      �?                      �?              �?                              $@              �?      @                      @              �?                      �?                       @               @       @      @                      @       @       @               @                               @              @      2@      7@      @      .@      7@              @      .@              @      @               @      @                      @               @       @               @                               @              @                               @      @      $@       @               @              @       @       @                      @      @       @      @      @       @      �?               @      �?              �?                      �?      �?              �?                              �?      @                                       @              @                      $@              �?      G@     �_@              7@      :@              7@      3@              5@      &@              @      @              @      @              @       @               @                      @       @              @      �?              �?      �?                      �?              �?                       @                              �?                      @                      �?              0@      @              ,@      @                       @              ,@      @              (@      �?              @                      @      �?              @                              �?               @       @                       @               @                       @                       @       @               @      @              �?                      �?      @                      @              �?      �?                      �?              �?                              @                      @      �?      7@     @Y@                      "@      �?      7@      W@      �?      .@     �@@      �?      *@      5@      �?      *@      3@      �?       @      3@              @      @                       @              @      �?                      �?              @              �?      @      0@              �?       @                      @              �?      @                      @              �?      �?                      �?              �?              �?      @       @               @      �?                      �?               @              �?       @      @               @              �?              @                      @      �?              �?      �?                                      �?              @                               @               @      (@                      (@               @                       @     �M@              @      I@                      3@              @      ?@               @      @                       @               @       @               @                               @              �?      ;@              �?      0@              �?                              0@                      &@              @      "@              @      @              @      @              �?                       @      @              �?      @              �?                              @              �?      �?              �?                              �?               @                              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�Bxg         �                   `_@^���?�           ��@       s                    �?20�����?�            �q@                           �?0����R�?_             b@                            �?r�q��?             8@������������������������       �                     @                          �U@��Q��?             4@������������������������       �                     �?                          pp@D�n�3�?             3@	                          P`@���!pc�?	             &@
                          �[@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           r@      �?              @������������������������       �                     @                          hr@      �?             @������������������������       �                      @                           \@      �?              @������������������������       �                     �?������������������������       �                     �?       `                    �?f�����?M             ^@       Q                    _@��n��d�??            @X@       *                   �_@����6�?6            @U@       )                   @^@-���?             ?@       (                   @q@:/����?             5@       !                   `\@�(\����?             4@                           �?��S�ۿ?	             .@������������������������       �                     "@                          `[@r�q��?             @������������������������       �                     @                           `Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @"       #                   @]@�Q����?             @������������������������       �                     �?$       '                   �U@      �?             @%       &                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@+       4                     �?����?!             K@,       3                   �d@�q�q�?             (@-       .                   �a@��(\���?             $@������������������������       �                     @/       2                   �c@�Q����?             @0       1                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @5       6                   �U@��g5��?             E@������������������������       �                      @7       B                   �e@��Q���?             D@8       A                   �a@������?	             ,@9       :                    `@VUUUUU�?             "@������������������������       �                     @;       @                    a@      �?             @<       ?                   @M@      �?             @=       >                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @C       J                   �c@�θ�?             :@D       E                   @l@�����H�?             2@������������������������       �                      @F       I                   �\@z�G�z�?             $@G       H                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @K       N                   �\@      �?              @L       M                   pd@���Q��?             @������������������������       �                      @������������������������       �                     @O       P                   �o@�q�q�?             @������������������������       �                      @������������������������       �                     �?R       S                   �Z@9��8���?	             (@������������������������       �                      @T       [                    �?ףp=
��?             $@U       Z                   @c@{�G�z�?             @V       W                   `k@      �?             @������������������������       �                     �?X       Y                   `@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?\       ]                   �a@z�G�z�?             @������������������������       �                     @^       _                   Pe@      �?              @������������������������       �                     �?������������������������       �                     �?a       h                   @[@�nkK�?             7@b       c                   �\@�$I�$I�?             @������������������������       �                      @d       e                     �?z�G�z�?             @������������������������       �                      @f       g                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?i       j                   �Y@      �?	             0@������������������������       �                     @k       r                    �?�q�q�?             (@l       m                     �?���|���?             &@������������������������       �                      @n       q                   �n@�<ݚ�?             "@o       p                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?t       }                     �?:���n�?Y            �a@u       |                   @|@�ʈD��?            �E@v       w                   @^@�(\����?             D@������������������������       �                    �@@x       y                   �d@؇���X�?             @������������������������       �                     @z       {                   �h@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @~       �                    @�TZa�?=            @X@       �                    �?��?"m�?7             U@�       �                   �]@8�Z$���?
             *@������������������������       �                     @�       �                   �a@h/�����?             "@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�Q����?             @�       �                   @e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   `@$JnY��?-            �Q@�       �                   �Z@���(\��?             $@������������������������       �                     @�       �                   �^@�$I�$I�?             @�       �                    �?�q�q�?             @�       �                   `\@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �^@H)h��8�?%            �N@�       �                    \@�U��nd�?              K@������������������������       �                     &@�       �                    �?G�6'�?            �E@�       �                    ]@d[����?            �B@������������������������       �                      @�       �                    �?Xnp�_��?            �A@�       �                   �]@      �?             @@������������������������       �                      @�       �                    �?R���Q�?             >@�       �                   �a@��JÝ�?             7@������������������������       �                     @�       �                   0e@�(\����?             4@�       �                   �d@�$I�$I�?             @�       �                   �c@z�G�z�?             @������������������������       �                     @�       �                   0k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     *@�       �                   b@؇���X�?             @������������������������       �                     @�       �                   d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �m@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �f@8�Z$���?             *@�       �                   `U@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                    `@��h�)�?(            |@�       �                    �?�P�n�?-             Q@������������������������       �                     @�       �                    �?�-ῃ�?(            �N@�       �                    �?p=
ףp�?             D@�       �                   �O@r�q��?             2@�       �                    `@@�0�!��?             1@�       �                   �Z@      �?             @������������������������       �                      @������������������������       �                      @�       �                    ^@$�q-�?             *@������������������������       �                     "@�       �                   P`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �_@j�V���?             6@������������������������       �                      @�       �                    �?z�G�z�?             4@�       �                   `]@X�<ݚ�?             "@������������������������       �                     @�       �                   �a@z�G�z�?             @������������������������       �                      @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                    �?�$I�$I�?             5@�       �                    �?p=
ףp�?             $@�       �                     �?r�q��?             @������������������������       �                      @�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @�       �                   `a@��!pc�?             &@�       �                    �?      �?             @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �?��]�b�?�            �w@�       o                  �a@��j�,��?�            `r@�                          �?
�H�h��?|            `f@�       �                   Pf@�*-x�!�?0            @Q@�       �                   �d@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�                         �c@     ��?-             P@�       �                    �?��ڊ�e�?%             I@�       �                   �[@$�q-�?	             *@������������������������       �                     �?������������������������       �                     (@�       �                   �S@��0\K5�?            �B@������������������������       �                     �?�                         �a@��ӭ�a�?             B@�       �                   Pa@H�7�&��?             >@�       �                    n@�����?             5@�       �                     �?"pc�
�?             &@�       �                    j@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        	             $@�                         �k@h/�����?             "@�                           ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        `]@r�q��?             @������������������������       �                     @                        �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        @`@      �?             @������������������������       �                     �?	      
                   a@���Q��?             @������������������������       �                      @                        (p@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          �?      �?             ,@������������������������       �                     �?                        �`@�	j*D�?             *@������������������������       �                     @                        0a@      �?              @������������������������       �                      @                        �d@�q�q�?             @������������������������       �                      @                        pe@      �?             @������������������������       �                      @������������������������       �                      @      6                    �?~��m�7�?L            �[@      1                  �p@h+�v:�?             A@      *                  pc@և���X�?             5@                         �?��
ц��?	             *@������������������������       �                     @      %                   �?���Q��?             $@      $                  @b@���Q��?             @       !                  �`@      �?             @������������������������       �                     �?"      #                  �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?&      '                  �]@���Q��?             @������������������������       �                      @(      )                  �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?+      ,                  pm@      �?              @������������������������       �                     @-      .                  �d@      �?             @������������������������       �                     �?/      0                  Pn@�q�q�?             @������������������������       �                      @������������������������       �                     �?2      3                   �?$�q-�?	             *@������������������������       �                     @4      5                   @r�q��?             @������������������������       �                     @������������������������       �                     �?7      J                   �?p���=�?5             S@8      A                  pc@�[��"e�?             2@9      <                   `@      �?             @:      ;                   �?      �?              @������������������������       �                     �?������������������������       �                     �?=      >                   �?      �?             @������������������������       �                     �??      @                  `b@�q�q�?             @������������������������       �                      @������������������������       �                     �?B      C                  �j@r�q��?	             (@������������������������       �                     @D      E                  0k@      �?              @������������������������       �                     �?F      G                  �p@؇���X�?             @������������������������       �                     @H      I                  pr@�q�q�?             @������������������������       �                     �?������������������������       �                      @K      L                  0`@^l��[B�?'             M@������������������������       �                     �?M      R                  @^@�MWl��?&            �L@N      Q                  `q@�q�q�?             @O      P                  @X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @S      l                  pf@@�0�!��?"            �I@T      U                  �l@�LQ�1	�?              G@������������������������       �                     5@V      ]                  �`@�+e�X�?             9@W      X                   b@؇���X�?             @������������������������       �                     @Y      Z                   �?      �?             @������������������������       �                     �?[      \                  @n@�q�q�?             @������������������������       �                     �?������������������������       �                      @^      _                  `n@�E��ӭ�?             2@������������������������       �                      @`      i                   @     ��?	             0@a      h                  �q@$�q-�?             *@b      g                   �?z�G�z�?             @c      d                  pa@�q�q�?             @������������������������       �                     �?e      f                  Pb@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @j      k                  q@�q�q�?             @������������������������       �                     �?������������������������       �                      @m      n                   @���Q��?             @������������������������       �                      @������������������������       �                     @p      �                   �?z.E���?F            �\@q      �                   �?he��#�?'            �N@r      s                   g@���]�`�?              J@������������������������       �                     @t      �                  �y@�?�K8��?            �H@u      z                   �?P���� �?             G@v      y                    �?z�G�z�?             $@w      x                  �c@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @{      �                  �d@0�����?             B@|      }                  c@�IєX�?             A@������������������������       �                     6@~                        (s@r�q��?	             (@������������������������       �                     @�      �                  `Z@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �                  �c@X�<ݚ�?             "@������������������������       �                      @�      �                  �c@����X�?             @�      �                  �m@r�q��?             @������������������������       �                     @�      �                  ``@�q�q�?             @�      �                  �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                  �j@���3L�?             K@������������������������       �                     (@�      �                   g@.0�w¹�?             E@�      �                  �l@�UH���?             C@�      �                   �?      �?              @������������������������       �                     @�      �                  �\@      �?             @�      �                  �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                   �?*;L]n�?             >@�      �                   �?`�Q��?             9@�      �                  �b@      �?              @������������������������       �                     @�      �                  @d@      �?             @������������������������       �                     @������������������������       �                     �?�      �                  @e@�t����?             1@�      �                   �?      �?             0@�      �                  p@�q�q�?             (@������������������������       �                      @�      �                  �a@z�G�z�?             $@������������������������       �                     @�      �                  �c@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                  0g@�|���?9             V@�      �                  �e@      �?             0@�      �                  �`@z�G�z�?             $@�      �                   e@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?      �?              @������������������������       �                     @�      �                  �b@z�G�z�?             @������������������������       �                      @�      �                  �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                   �?~X�<��?.             R@�      �                  0b@b-�I�w�?             C@�      �                  pb@��Θ���?             =@�      �                  �i@�K8��?             :@�      �                   `@      �?             @������������������������       �                     �?�      �                  `@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  0l@���7�?             6@�      �                   `@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@������������������������       �                     @�      �                  �d@h/�����?             "@������������������������       �                     @�      �                  i@VUUUUU�?             @������������������������       �                      @�      �                  �q@      �?             @������������������������       �                      @������������������������       �                      @�      �                  �`@г�wY;�?             A@������������������������       �                     =@�      �                  �i@z�G�z�?             @������������������������       �                     @�      �                  @b@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KM�KK��h[�BX,       �J@     �v@      t@      =@      \@     �a@      6@     @R@     �H@      �?       @      .@                      @      �?       @      &@      �?                               @      &@              @       @              @      �?                      �?              @                              @              @      @              @                      �?      @                       @              �?      �?              �?                              �?      5@     @P@      A@      1@      L@      8@      *@     �J@      3@       @      ;@       @       @      1@       @      �?      1@       @              ,@      �?              "@                      @      �?              @                       @      �?                      �?               @              �?      @      �?      �?                              @      �?               @      �?               @                              �?              �?              �?                              $@              &@      :@      1@      �?      @       @      �?      �?       @                      @      �?      �?      @      �?      �?                      �?              �?                                      @               @              $@      7@      "@       @                       @      7@      "@       @      @      @      @      @      @      @                              @      @              @      �?              �?      �?                      �?              �?                       @                               @      @                              4@      @              0@       @               @                       @       @              �?       @                       @              �?                      @                      @      @              @       @                       @              @                      �?       @                       @              �?              @      @      @       @                       @      @      @       @       @      �?       @       @                      �?               @      �?                      �?               @                                      �?              �?      @                      @              �?      �?              �?                              �?      @      "@      $@      @      �?       @                       @      @      �?               @                       @      �?               @                              �?                       @       @                      @               @      @              @      @                       @              @       @              �?       @              �?                               @              @                      �?              @     �C@     �W@              @     �C@              �?     �C@                     �@@              �?      @                      @              �?       @                       @              �?                      @              @     �A@     �K@      @      8@     �J@      �?       @      @              @              �?      @      @              �?      @              �?                              @      �?      @      �?              @      �?              @                              �?      �?                      @      0@     �H@      @      @      �?              @              @       @      �?      @       @               @      �?                      �?               @                       @      �?               @                              �?                              �?       @      &@      H@       @      @     �F@                      &@       @      @      A@       @      @      <@               @               @      @      <@       @      @      9@                       @       @      @      7@       @      @      1@              @               @      �?      1@       @      �?      @              �?      @                      @              �?      �?                      �?              �?               @                                      *@              �?      @                      @              �?       @              �?                               @                      @                      @              @      @              @                              @              &@       @              �?       @              �?                               @              $@              8@      o@      f@      @     �H@      .@              @              @      E@      .@       @      ?@      @              .@      @              ,@      @               @       @               @                               @              (@      �?              "@                      @      �?                      �?              @                      �?               @      0@      @       @                              0@      @              @      @              @                      �?      @                       @              �?       @              �?                               @              &@               @      &@       @      �?       @      @      �?              @                       @      �?              @      �?                                      @               @       @               @                               @      �?      "@      �?      �?       @      �?      �?              �?      �?                                      �?               @                      @              4@      i@     @d@      1@     �a@      a@      @      S@     @X@      @      F@      4@              �?      @              �?                              @      @     �E@      0@      @     �C@      @      �?      (@              �?                              (@              @      ;@      @      �?                       @      ;@      @       @      8@      @              3@       @              "@       @              �?       @              �?                               @               @                      $@               @      @       @       @              �?       @                                      �?              @      �?              @                       @      �?                      �?               @                      @      @              �?                       @      @                       @               @      �?                      �?               @              �?      @      "@      �?                              @      "@                      @              @      @               @                       @      @                       @               @       @               @                               @      �?      @@     @S@              *@      5@              (@      "@              @      @                      @              @      @              @       @              @      �?              �?                       @      �?                      �?               @                              �?              @       @               @                      �?       @                       @              �?                      @       @              @                       @       @              �?                      �?       @                       @              �?                      �?      (@                      @              �?      @                      @              �?              �?      3@      L@      �?      @      &@      �?      @      �?              �?      �?              �?                              �?      �?      @                      �?              �?       @                       @              �?                               @      $@                      @               @      @              �?                      �?      @                      @              �?       @              �?                               @              *@     �F@                      �?              *@      F@              @       @              �?       @              �?                               @              @                      "@      E@              @      D@                      5@              @      3@              �?      @                      @              �?      @                      �?              �?       @              �?                               @              @      *@               @                      @      *@              �?      (@              �?      @              �?       @                      �?              �?      �?              �?                              �?                       @                       @               @      �?                      �?               @                      @       @                       @              @              &@      P@      D@      $@      F@      @      @      D@      @      @                       @      D@      @       @      D@      @               @       @              @       @              @                               @              @               @      @@       @       @      @@                      6@               @      $@                      @               @      @                      @               @                                       @                      @      @      @                       @              @       @              @      �?              @                       @      �?              �?      �?              �?                              �?              �?                              �?              �?      4@     �@@                      (@      �?      4@      5@      �?      4@      1@      �?      @                      @              �?      @              �?      �?                      �?              �?                               @                      *@      1@               @      1@              @      @                      @              @      �?              @                              �?              @      (@              @      (@              @       @               @                       @       @                      @               @      @               @                              @                      @              �?                      @                              @      @      N@      9@               @      ,@               @       @              �?      �?                      �?              �?                      �?      @                      @              �?      @                       @              �?       @              �?                               @                      @      @      M@      &@      @      9@      $@      �?      7@      @      �?      7@       @               @       @              �?                      �?       @              �?                               @      �?      5@              �?      @              �?                              @                      ,@                              @       @       @      @                      @       @       @       @       @                               @       @                       @               @                     �@@      �?              =@                      @      �?              @                      �?      �?                      �?              �?        �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJQY%hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�i         �                   �c@�����?�           ��@       C                   `_@.1���?i            �c@       B                    W@\Ư�,�?/            @Q@       	                     �?     ��?,             P@                          �Y@�q�q�?             @������������������������       �                      @                           �?      �?             @������������������������       �                      @������������������������       �                      @
       %                   `]@R[4�0`�?)             M@                          �`@�ങa�?             ?@                           \@��JÝ�?             7@                           �?{�G�z�?             @������������������������       �                      @                          �Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          @^@r�q��?             2@������������������������       �                     "@                          �^@�q�q�?             "@������������������������       �                     �?                          �_@      �?              @������������������������       �                      @                          P`@�q�q�?             @                          �[@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                     �?       $                    �?      �?              @       !                    �?������?             @                           @Z@      �?             @������������������������       �                     @������������������������       �                     �?"       #                   Pb@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?&       )                    �?�n���?             ;@'       (                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?*       =                   �c@�8��8��?             8@+       :                   �^@R��Xp�?             3@,       9                   @^@
ц�s�?
             *@-       4                    �?�8��8��?	             (@.       3                   �[@      �?              @/       2                    �?      �?             @0       1                    X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @5       8                    �?      �?             @6       7                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?;       <                   �Z@r�q��?             @������������������������       �                     �?������������������������       �                     @>       A                    �?z�G�z�?             @?       @                   Pe@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @D       {                   Pc@|CX�D��?:            @V@E       h                    �?2�tk~X�?0             R@F       g                   �d@FGr���?!             I@G       T                   �`@�q�q��?              H@H       M                    `@�E�_���?             5@I       J                   �_@z�G�z�?             @������������������������       �                     �?K       L                    ]@      �?             @������������������������       �                     �?������������������������       �                     @N       O                    �?      �?             0@������������������������       �                     $@P       Q                   �^@r�q��?             @������������������������       �                     @R       S                   Pb@      �?              @������������������������       �                     �?������������������������       �                     �?U       `                    �?l��
I��?             ;@V       _                   �a@"pc�
�?	             &@W       ^                   `Q@      �?              @X       Y                   `R@�q�q�?             @������������������������       �                     �?Z       [                    �?z�G�z�?             @������������������������       �                     @\       ]                   0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @a       f                    �?      �?             0@b       c                    a@�q�q�?             "@������������������������       �                     @d       e                    _@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @i       z                   �a@�J����?             6@j       y                    I@0\�Uo��?             3@k       x                    @     ��?             0@l       q                    �?�q-��?	             *@m       p                   �]@�Q����?             @n       o                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r       u                   �]@      �?              @s       t                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @v       w                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @|       }                    �?�IєX�?
             1@������������������������       �                      @~       �                   �^@�����H�?             "@       �                     �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       6                   �?�"e��b�?r            �@�       �                     �?�v����?�            r@�       �                    �?$߼�x�?!             N@�       �                   �`@N���-��?             �M@�       �                   �^@П[;U��?             =@�       �                    \@      �?              @������������������������       �                     @�       �                   @b@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �a@�q�q�?	             5@�       �                   �k@�<ݚ�?             "@������������������������       �                     @�       �                   @Z@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     (@�       �                    c@�d��0�?             >@�       �                   �g@P���Q�?             4@������������������������       �                     �?������������������������       �                     3@�       �                   xv@      �?             $@�       �                   pc@����X�?             @�       �                   �q@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       )                  0c@lċ��?�            �l@�       (                  �}@�n>.L!�?�            `i@�       #                  �u@$��7e�?            �h@�                          �?�R��J��?z            �g@�       �                    a@���s���?j            �d@�       �                   @Z@�W��#V�?<             W@������������������������       �                      @�       �                    �?F@����?:            �V@�       �                   �q@��^B{	�?/             R@�       �                    �?�5	h�c�?+            @P@�       �                    j@<�
I��?             3@������������������������       �                     @�       �                   @^@0�����?             ,@�       �                   `k@      �?             @������������������������       �                     �?�       �                   �Z@�q�q�?             @������������������������       �                     �?�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `\@ףp=
�?             $@�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �`@P���� �?             G@�       �                    _@ ��WV�?             :@������������������������       �        	             .@�       �                   �k@�C��2(�?             &@������������������������       �                     @�       �                   �_@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �\@�Q����?             4@�       �                   �[@�q�q�?             "@�       �                   Hp@؇���X�?             @������������������������       �                     @�       �                   �W@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   �^@"pc�
�?             &@������������������������       �                     @�       �                   �k@����X�?             @������������������������       �                      @������������������������       �                     @�       �                   �^@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �^@r�q��?             2@�       �                   �V@      �?             @������������������������       �                      @������������������������       �                      @�       �                    _@@4և���?	             ,@������������������������       �                     &@�       �                   �g@�q�q�?             @������������������������       �                     �?�       �                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   Pc@���^B{�?.             R@�       �                   pf@6M5���?            �D@�       �                    �?r�q��?             @�       �                   �e@z�G�z�?             @�       �                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �b@<=�,S��?            �A@�       �                    �?��
ц��?             :@������������������������       �                     @�       �                   �[@և���X�?             5@�       �                   �a@����X�?             @�       �                   �m@�q�q�?             @������������������������       �                     @�       �                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �a@����X�?	             ,@�       �                    �?      �?              @�       �                   Hp@և���X�?             @������������������������       �                     @�       �                   @_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �b@�����H�?             "@������������������������       �                     @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?                          e@�n`���?             ?@                         �?�IєX�?             1@������������������������       �                     @                         d@�8��8��?             (@������������������������       �                     @      
                  0d@      �?              @                        p`@z�G�z�?             @������������������������       �                      @      	                  �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                        �^@X�Cc�?             ,@������������������������       �                     @                        Pe@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@                         �?�g\��?             :@                         �?@�0�!��?             1@                        �r@r�q��?             @������������������������       �                     @������������������������       �                     �?                        �]@"pc�
�?             &@������������������������       �                     @                        Pk@���Q��?             @������������������������       �                      @                        �^@�q�q�?             @������������������������       �                     �?                        pq@      �?              @������������������������       �                     �?������������������������       �                     �?                          `@�<ݚ�?             "@������������������������       �                     @!      "                  �k@�q�q�?             @������������������������       �                     �?������������������������       �                      @$      '                  0{@0�����?             @%      &                   `@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @*      5                  `t@�θ�?             :@+      0                  �[@�z�G��?             4@,      /                   g@$�q-�?	             *@-      .                  �U@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@1      2                  �d@����X�?             @������������������������       �                     @3      4                  �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @7      ^                   _@Oo�f��?�            �q@8      W                   �?\�5��?#             J@9      P                   b@z�5���?             C@:      I                  0q@X�<ݚ�?             ;@;      @                  �j@�E��ӭ�?             2@<      =                   �?z�G�z�?             @������������������������       �                      @>      ?                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?A      H                   �?$�q-�?             *@B      G                  @`@�����H�?             "@C      F                   �?z�G�z�?             @D      E                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @J      O                   �?�<ݚ�?             "@K      N                    �?      �?              @L      M                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?Q      V                  �o@���k���?             &@R      U                    �?�<ݚ�?             "@S      T                  `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @X      ]                   @����S�?
             ,@Y      \                  @]@$�q-�?	             *@Z      [                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     �?_      �                  0e@�m��G-�?�            `m@`      �                   �?61m#�?v             g@a      n                  �o@t����{�?            �B@b      k                   �?�IєX�?             1@c      f                   �?؇���X�?	             ,@d      e                  pm@      �?              @������������������������       �                     �?������������������������       �                     �?g      j                   @�8��8��?             (@h      i                   b@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @l      m                  �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @o      p                  �`@{�G�z�?             4@������������������������       �                     @q      �                  hr@     ��?             0@r      w                  8q@*D>��?
             *@s      t                  �_@�Q����?             @������������������������       �                     �?u      v                  0b@      �?             @������������������������       �                     �?������������������������       �                     @x      y                  �q@      �?              @������������������������       �                      @z                         d@�q�q�?             @{      ~                    �?z�G�z�?             @|      }                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                  �`@D˩�m��?]            �b@�      �                   @Rԅ5l�?A            @[@�      �                   �?��Dl<�?>            �Z@�      �                   q@@S�)�q�?6            �V@�      �                   d@���L��?-            �Q@�      �                   `@     ��?*             P@�      �                  �p@"Ae���?            �G@�      �                   �?^����?            �E@�      �                   �?��a�n`�?             ?@�      �                  �j@R�}e�.�?             :@�      �                  �g@ףp=
�?	             $@�      �                  �f@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                    �?      �?             0@������������������������       �                     �?�      �                  �^@���Q��?             .@�      �                  �\@z�G�z�?             @������������������������       �                     �?�      �                  �o@      �?             @������������������������       �                     �?������������������������       �                     @�      �                  �a@z�G�z�?             $@������������������������       �                     @�      �                  �m@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�      �                  0k@�q�q�?             (@�      �                  �g@r�q��?             @������������������������       �                     �?������������������������       �                     @�      �                    �?�q�q�?             @������������������������       �                     �?�      �                  �b@���Q��?             @������������������������       �                      @�      �                  �\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   �?�IєX�?             1@������������������������       �                     @�      �                  pb@@4և���?	             ,@�      �                    �?z�G�z�?             @�      �                  �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     @������������������������       �        	             5@������������������������       �                     .@�      �                  �_@�q�q�?             @������������������������       �                     �?�      �                  0c@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?�n_Y�K�?            �C@�      �                  �`@���B���?             :@������������������������       �                     �?�      �                   `@�J�4�?             9@������������������������       �                     �?�      �                  Pb@      �?             8@�      �                  `c@���!pc�?             &@�      �                  �k@      �?              @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                  a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             *@�      �                   r@�θ�?	             *@�      �                  @a@�C��2(�?             &@������������������������       �                     @�      �                   b@      �?              @�      �                  �b@z�G�z�?             @������������������������       �                      @�      �                  0d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�      �                  �n@���QI�?$             I@������������������������       �                     <@�      �                  `o@�0�~�4�?             6@������������������������       �                     �?�      �                   @�����?             5@�      �                  �e@P���Q�?             4@������������������������       �        	             &@�      �                   q@�����H�?             "@�      �                  �^@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KM�KK��h[�BH-        I@     �v@     �s@      7@     �X@      B@      1@      A@      2@      1@      =@      2@      @       @               @                       @       @                       @               @                      *@      ;@      2@      @      2@      @      @      1@       @      �?       @       @               @              �?               @      �?                                       @      @      .@                      "@              @      @              �?                       @      @                       @               @      @               @      @              �?                      �?      @                      �?              @      �?      @      @      �?      @      @              �?      @                                      �?              �?       @                       @              �?                              �?      @      "@      (@       @      �?               @                              �?              @       @      (@      @      @      &@      @      @      @       @      @      @      �?      �?      @      �?      �?       @      �?               @                       @      �?                              �?                              @      �?      @              �?       @                       @              �?                              �?              �?                      �?              @      �?                                      @              @      �?              @      �?              @                              �?              �?                      @              @     @P@      2@      @     �H@      1@      �?      C@      &@      �?      C@      "@      �?      3@      �?              @      �?              �?                      @      �?                      �?              @              �?      .@                      $@              �?      @                      @              �?      �?              �?                              �?                      3@       @              "@       @              @       @              @       @                      �?              @      �?              @                      �?      �?              �?                              �?               @                      @                      $@      @              @      @                      @              @      @              @                              @              @                               @      @      &@      @      @       @      @      @       @      @      @      @      @      @      �?      �?              �?      �?                      �?              �?              @                       @      @       @       @      �?                      �?               @                              @       @                       @              @                      @                              @              @                      0@      �?               @                       @      �?              @      �?                      �?              @                      @              ;@     �p@     �q@      5@     `g@     @T@      �?      C@      5@      �?     �B@      5@              *@      0@              @       @              @                      �?       @                       @              �?                      @      ,@              @       @              @                       @       @                       @               @                              (@      �?      8@      @      �?      3@              �?                              3@                      @      @               @      @              �?      @              �?                              @              �?      �?                      �?              �?                      @                      �?              4@     �b@      N@      ,@      `@      N@      ,@     �^@      N@      *@     �^@     �K@      &@     @Y@      J@      $@     @R@      "@                       @      $@     @R@      @      $@      M@      @      @     �K@      @       @      .@       @              @               @      $@       @       @      �?      �?                      �?       @      �?              �?                      �?      �?                      �?              �?                              "@      �?              �?      �?              �?                              �?               @              @      D@       @      �?      9@                      .@              �?      $@                      @              �?      @              �?                              @              @      .@       @      @      @              �?      @                      @              �?       @                       @              �?                       @                              "@       @              @                      @       @                       @              @              @      @              @                              @                      .@      @               @       @                       @               @                      *@      �?              &@                       @      �?              �?                      �?      �?                      �?              �?              �?      <@     �E@      �?      6@      2@      �?              @      �?              @      �?               @      �?                                       @                       @                      �?              6@      *@              ,@      (@              @                      "@      (@              @       @              @       @              @                      �?       @                       @              �?                      �?                      @      $@              @      @              @      @              @                      �?      @                      @              �?                              �?                      @               @      �?              @                      �?      �?              �?                              �?              @      9@              �?      0@                      @              �?      &@                      @              �?      @              �?      @                       @              �?       @              �?                               @                      @              @      "@              @                       @      "@               @                              "@       @      5@      @              ,@      @              @      �?              @                              �?              "@       @              @                      @       @               @                      �?       @                      �?              �?      �?                      �?              �?               @      @                      @               @      �?                      �?               @                      �?      �?      @              �?      @              �?                              @      �?                              @              @      4@              @      ,@              �?      (@              �?       @              �?                               @                      $@              @       @              @                       @       @                       @               @                              @              @     @T@      i@      @      :@      7@       @      ,@      6@              (@      .@              @      *@              @      �?               @                       @      �?               @                              �?              �?      (@              �?       @              �?      @              �?      @                      @              �?                              �?                      @                      @              @       @              @      �?              �?      �?                      �?              �?                      @                              �?       @       @      @       @              @       @              �?       @                                      �?                      @               @              �?      (@      �?              (@      �?               @      �?                      �?               @                      $@              �?                      @     �K@      f@       @     �J@     @`@       @      3@      0@      �?      (@      @              (@       @              �?      �?                      �?              �?                      &@      �?               @      �?               @                              �?              @              �?               @      �?                                       @      �?      @      (@                      @      �?      @       @      �?      @      @      �?      �?      @      �?                              �?      @              �?                              @              @       @               @                      @       @              @      �?              �?      �?              �?                              �?              @                              �?                      @              A@     �\@              3@     �V@              1@     @V@              1@     �R@              1@     �J@              1@     �G@              0@      ?@              (@      ?@              @      8@              @      3@              �?      "@              �?      @                      @              �?                              @              @      $@                      �?              @      "@              @      �?              �?                      @      �?                      �?              @                       @       @                      @               @      @               @                              @                      @              @      @              �?      @              �?                              @              @       @              �?                      @       @               @                      �?       @                       @              �?                      @                      �?      0@                      @              �?      *@              �?      @              �?       @                       @              �?                               @                      "@                      @                      5@                      .@               @      �?              �?                      �?      �?              �?                              �?              .@      8@              @      5@              �?                      @      5@              �?                      @      5@              @       @              �?      @              �?      �?              �?                              �?                      @               @      �?                      �?               @                              *@              $@      @              $@      �?              @                      @      �?              @      �?               @                       @      �?                      �?               @                      @                               @      �?       @     �G@                      <@      �?       @      3@      �?                               @      3@              �?      3@                      &@              �?       @              �?      @              �?                              @                      @              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��fbhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�l         �                   �`@z+`�K�?�           ��@       �                    �?���Bk�?�            �r@       b                    �?V;�����?�             l@       %                   �h@�>��*�?d            �b@                            �?t��*f��?             E@������������������������       �                     @       "                   �b@��Ha���?            �C@       !                   �g@pB躍�?             A@	       
                   �Y@     ��?             @@������������������������       �                     @                          g@��1+��?             ;@                          `[@�^)��?             9@                          �_@      �?             @������������������������       �                      @                          @`@      �?              @������������������������       �                     �?������������������������       �                     �?                          �e@0�����?             5@                          �]@�)O�?             2@������������������������       �                     @                           `@�g���e�?             &@                           �?������?             @                          �]@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                          �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @#       $                   �V@z�G�z�?             @������������������������       �                     �?������������������������       �                     @&       7                    �?!r�i��?E             [@'       (                   �Y@r�q��?             8@������������������������       �                     @)       ,                    \@p=
ףp�?             4@*       +                   �a@���Q��?             @������������������������       �                     @������������������������       �                      @-       2                   p`@���Q��?             .@.       1                   pl@�8��8��?             (@/       0                    _@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @3       4                    j@�q�q�?             @������������������������       �                     �?5       6                   `@      �?              @������������������������       �                     �?������������������������       �                     �?8       O                    �?��8��8�?6             U@9       L                   c@P��)x9�?'             L@:       ;                     �?���QI�?#             I@������������������������       �                     @<       G                   �k@0'�%���?              G@=       @                   �Y@      �?             0@>       ?                   p`@�q�q�?             @������������������������       �                      @������������������������       �                     �?A       F                    ]@$�q-�?	             *@B       E                   �a@r�q��?             @C       D                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @H       K                   �\@(;L]n�?             >@I       J                   �\@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     :@M       N                   �c@r�q��?             @������������������������       �                     �?������������������������       �                     @P       a                   `^@h�����?             <@Q       X                   �]@և���X�?             5@R       S                     �?�����H�?             "@������������������������       �                     @T       W                   �V@r�q��?             @U       V                    U@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @Y       \                   �q@�8��8��?             (@Z       [                   po@���Q��?             @������������������������       �                      @������������������������       �                     @]       ^                     �?؇���X�?             @������������������������       �                      @_       `                   pr@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @c       �                   �_@ʝ]o9"�?1            �R@d                          �^@˒���G�?             C@e       ~                   Hp@.�?�P��?             >@f       o                   �[@�-Z0�?             =@g       n                   @]@�h$��W�?             .@h       m                   `[@�Q����?             $@i       l                    [@{�G�z�?             @j       k                    `@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @p       }                    �?/����?	             ,@q       r                    Y@�θ�?             *@������������������������       �                     @s       |                    `@�z�G��?             $@t       u                   �Z@և���X�?             @������������������������       �                     �?v       w                   `\@�q�q�?             @������������������������       �                     �?x       {                    \@���Q��?             @y       z                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    ^@:Mw;�?            �B@�       �                   @c@�nkK�?             7@������������������������       �        
             .@�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     @�       �                   Pa@*x9/��?             ,@������������������������       �                     @�       �                   �^@      �?              @������������������������       �                      @�       �                   pm@�8��8��?             @������������������������       �                     @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @Z@(�@݈g�?6             S@������������������������       �                     @�       �                   �]@��_�Qv�?4            @R@�       �                   �]@|L�Sw�?            �A@�       �                   @]@����e��?            �@@�       �                    �?     ��?             @@�       �                   0a@      �?             8@�       �                   �Z@���ĳ��?             .@�       �                     �?���|���?
             &@�       �                   @X@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @Y@�q�q�?             "@�       �                   @\@և���X�?             @������������������������       �                     �?�       �                   @_@�q�q�?             @�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                     �?      �?             @�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�����H�?             "@������������������������       �                      @�       �                   �i@؇���X�?             @�       �                   �W@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   ``@z�5���?             C@�       �                     �?dG�+�?             ?@������������������������       �                      @�       �                   �a@h�d0ܩ�?             7@�       �                    �?�8��8��?	             (@�       �                    [@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �Q@      �?              @�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �c@      �?             @������������������������       �                     �?�       �                    �?���Q��?             @�       �                   `^@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    _@"pc�
�?             &@�       �                    �?����X�?             @������������������������       �                     @�       �                   `X@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?؇���X�?             @�       �                   �_@r�q��?             @�       �                   �\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                  �c@�W��p�?           {@�       �                  0e@z_R��:�?�            �x@�                          �?�s��:��?�             s@�       �                     �?V�dD��?)            �M@�       �                   Pg@&�'+�>�?             ?@������������������������       �                     @�       �                    @�:����?             ;@�       �                   �`@g\�5�?             :@�       �                   �c@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�       �                   �m@���ĳ��?             .@�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   q@j�V���?	             &@�       �                   pp@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    b@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   @i@������?             <@�       �                   �\@�8��8��?             @������������������������       �                     �?�       �                   `h@���Q��?             @������������������������       �                      @������������������������       �                     @�                          @�i�V��?             6@�       �                   0l@6�����?             5@������������������������       �                     @�       �                   Pa@�M�]��?             1@������������������������       �                      @�                          �a@���ĳ��?             .@������������������������       �                      @                        0c@&�q-�?             *@                        �]@�Q����?             @������������������������       �                      @                         b@VUUUUU�?             @������������������������       �                     �?                        �b@      �?              @������������������������       �                     �?������������������������       �                     �?	                        `r@      �?              @
                        Pp@����X�?             @                        �c@���Q��?             @������������������������       �                     �?                        �[@      �?             @������������������������       �                     �?                        �l@�q�q�?             @������������������������       �                     �?                        �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?      4                   I@$��N���?�            �n@      +                   �?���(\��?             >@      *                  �^@��[r��?             5@                        `X@9��8���?	             (@                         �?      �?             @������������������������       �                     �?                        b@�q�q�?             @������������������������       �                     �?������������������������       �                      @       %                   c@      �?              @!      "                   �?      �?             @������������������������       �                     �?#      $                  �[@�q�q�?             @������������������������       �                     �?������������������������       �                      @&      '                  �Z@      �?             @������������������������       �                     �?(      )                   \@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@,      /                   �?X�<ݚ�?             "@-      .                   �?      �?             @������������������������       �                     �?������������������������       �                     @0      3                   �?���Q��?             @1      2                   @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?5      @                  �f@��ò���?�            �j@6      ?                   �?T���N@�?             9@7      8                  �`@�������?             (@������������������������       �                     �?9      :                  �d@�C��2(�?             &@������������������������       �                     @;      <                  �a@r�q��?             @������������������������       �                     @=      >                   c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             *@A      �                  �d@ư���?�?r            �g@B      �                   �?Rj��	��?m            �f@C      x                   �?
ףp=
�?c             d@D      s                   �?-a���?+            �P@E      j                  Pc@������?$            �M@F      M                  �j@ȩm��?            �F@G      H                  0b@���|���?             &@������������������������       �                     @I      J                  @_@z�G�z�?             @������������������������       �                      @K      L                  `g@�q�q�?             @������������������������       �                     �?������������������������       �                      @N      W                   o@�M�]��?             A@O      P                  0a@      �?	             ,@������������������������       �                     �?Q      T                    �?�؉�؉�?             *@R      S                  @b@      �?             @������������������������       �                     �?������������������������       �                     @U      V                  �a@�q�q�?             "@������������������������       �                     @������������������������       �                     @X      Y                  `p@�G�z��?             4@������������������������       �                     @Z      [                  �p@ҳ�wY;�?             1@������������������������       �                     @\      g                  ``@և���X�?	             ,@]      `                  0q@�z�G��?             $@^      _                  Pb@�q�q�?             @������������������������       �                      @������������������������       �                     �?a      b                   ^@؇���X�?             @������������������������       �                      @c      f                  �a@z�G�z�?             @d      e                  8s@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @h      i                  �q@      �?             @������������������������       �                     �?������������������������       �                     @k      l                  �h@����X�?	             ,@������������������������       �                      @m      n                    �?r�q��?             (@������������������������       �                     @o      p                  �k@�<ݚ�?             "@������������������������       �                     @q      r                  d@���Q��?             @������������������������       �                     @������������������������       �                      @t      w                  Pb@      �?              @u      v                   b@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @y      �                  pd@�חF�P�?8            @W@z      {                  �j@�k��?6            @V@������������������������       �                     4@|      �                  �m@��X���?+            @Q@}      �                   �?�LQ�1	�?             7@~                         �?�q�q�?             5@������������������������       �                     @�      �                  �[@��S���?	             .@������������������������       �                     @�      �                   @���|���?             &@�      �                  �a@���Q��?             $@������������������������       �                      @�      �                  �c@      �?              @�      �                  @_@؇���X�?             @�      �                  �l@r�q��?             @������������������������       �                     @�      �                  0m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                  �\@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  �`@�q��/��?             G@�      �                  �^@г�wY;�?             A@�      �                   q@���N8�?             5@�      �                   �?؇���X�?             @�      �                    �?r�q��?             @������������������������       �                     �?�      �                  �\@z�G�z�?             @������������������������       �                     �?�      �                  �o@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@������������������������       �                     *@�      �                   @�q�q�?
             (@�      �                    �?      �?              @�      �                  0a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �                  q@      �?             @������������������������       �                      @������������������������       �                      @�      �                  ``@      �?             @������������������������       �                      @������������������������       �                      @�      �                  �^@�G�z��?
             4@������������������������       �                     @�      �                  0c@     ��?             0@�      �                  �r@      �?              @�      �                   �?r�q��?             @������������������������       �                     �?�      �                  �m@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                   �?      �?              @������������������������       �                     @������������������������       �                      @�      �                  pl@H�z�G�?             $@������������������������       �                     @�      �                   o@      �?             @������������������������       �                     @������������������������       �                     �?�      �                  �c@pY�^;�?8            �W@�      �                   �?��Kh/�?	             2@�      �                  �[@      �?              @������������������������       �                      @������������������������       �                     @�      �                  �`@      �?             $@�      �                   �?r�q��?             @������������������������       �                      @�      �                  �O@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                  Hq@��}���?/            @S@�      �                  a@�>����?#             K@�      �                  �`@ףp=
�?             D@�      �                  �i@�L���?            �B@������������������������       �                     *@�      �                   �?      �?             8@������������������������       �                      @�      �                    �?��2(&�?             6@�      �                   �?      �?             @������������������������       �                     �?�      �                  pe@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?�X�<ݺ?
             2@�      �                  n@      �?             0@������������������������       �                     "@�      �                   �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                  `e@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             ,@�      �                  `r@��+7��?             7@�      �                   �?z�G�z�?             @������������������������       �                      @�      �                  `e@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                  �f@�����H�?	             2@������������������������       �                     0@������������������������       �                      @�      �                  d@��wY;�?             A@�      �                   �?PN��T'�?             ;@�      �                   �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �        	             3@������������������������       �                     @�t�b�      h�h(h+K ��h-��R�(KM�KK��h[�B�.        N@     u@     u@      ?@      i@     @Q@      8@     `d@      C@      0@     �\@      4@      @      9@      &@              @              @      6@      &@      @      6@      @      @      6@      @              @              @      1@      @      @      0@      @       @      �?      �?       @                              �?      �?                      �?              �?              @      .@      @      �?      ,@      @              @              �?      @      @      �?      @      @              @      @              @                              @      �?                              @               @      �?                      �?               @                              �?      �?              �?                              �?                       @      �?              @      �?                                      @      $@     @V@      "@      @      0@      @      @                      �?      0@      @              @       @              @                               @      �?      *@      �?      �?      &@              �?      @              �?                              @                      @                       @      �?              �?                      �?      �?                      �?              �?              @     @R@      @      @      J@      �?       @     �G@      �?              @               @     �E@      �?      �?      ,@      �?               @      �?               @                              �?      �?      (@              �?      @              �?       @                       @              �?                              @                      @              �?      =@              �?      @              �?                              @                      :@              �?      @              �?                              @               @      5@      @       @      ,@      @               @      �?              @                      @      �?              �?      �?              �?                              �?              @               @      @      @       @              @       @                                      @              @      �?               @                      @      �?              @                              �?              @               @     �H@      2@      @      2@      .@      @      2@      @      @      1@      @       @      @      @       @       @      @       @       @      �?       @              �?       @                                      �?               @                              @              @              @      $@      �?      @      $@                      @              @      @              @      @              �?                       @      @                      �?               @      @              �?       @              �?                               @              �?      �?                      @                              �?              �?                               @      @      ?@      @      �?      6@                      .@              �?      @              �?                              @               @      "@      @              @               @      @      @                       @       @      @      �?              @               @              �?                      �?       @                      @      C@      ?@      @                      @      C@      ?@       @      8@      "@       @      6@      "@       @      6@       @      �?      0@      @      �?       @      @              @      @              �?      �?                      �?              �?                      @      @              @      @                      �?              @       @              @      �?               @                       @      �?               @                              �?                      �?               @              �?      �?       @              �?      �?              �?                              �?      �?              �?                      �?      �?                               @      �?               @                      @      �?              �?      �?              �?                              �?              @              �?      @      �?              @              �?              �?                      �?      �?                                      �?               @               @      ,@      6@       @       @      5@                       @       @       @      *@       @      @      @      �?      @              �?                              @              �?      @      @      �?              �?                      �?      �?                              @      @              �?                       @      @              �?      @              �?                              @              �?                       @      "@               @      @                      @               @       @               @                               @                      @              @      �?              @      �?               @      �?               @                              �?              @                      �?              =@      a@     �p@      9@     @\@     Pp@      7@     �X@     �f@      $@      6@      ;@      @      &@      ,@      @                       @      &@      ,@       @      &@      *@               @      "@                      "@               @               @      "@      @              �?      @                      @              �?               @       @      �?       @      @                      @               @                              @      �?                      �?              @                              �?      @      &@      *@      @       @      �?                      �?      @       @                       @              @                      �?      "@      (@      �?       @      (@                      @      �?       @       @                       @      �?       @      @               @              �?      @      @      �?      �?      @                       @      �?      �?      �?                      �?      �?      �?                      �?              �?                              @      @              @       @              @       @              �?                       @       @                      �?               @      �?              �?                      �?      �?              �?                              �?               @                              �?              �?              *@      S@     �c@      @      1@       @      @      (@      @      @      @      @      @              �?      �?                       @              �?                      �?       @                       @      @      @       @      �?      �?                      �?       @      �?                      �?               @                               @       @                      �?               @      �?               @                              �?              "@                      @      @              @      �?                      �?              @                       @      @              �?      @                      @              �?                      �?               @     �M@     �b@      �?      �?      7@      �?      �?      $@              �?              �?              $@                      @      �?              @                      @      �?              �?      �?                                      �?                      *@      @      M@     @_@      @     �L@     �]@      @      H@      [@      @     �@@      >@      @      <@      ;@      @      8@      1@              @      @                      @              @      �?               @                       @      �?                      �?               @              @      4@      $@      @      "@      �?      �?                      @      "@      �?              @      �?                      �?              @              @      @                      @              @                              &@      "@                      @              &@      @              @                       @      @              @      @              �?       @                       @              �?                      @      �?               @                      @      �?              �?      �?                      �?              �?                      @                      �?      @              �?                              @              @      $@               @                       @      $@                      @               @      @                      @               @      @                      @               @                      @      @              @      �?              @                              �?                       @              .@     �S@              *@      S@                      4@              *@      L@               @      .@              @      ,@                      @              @       @                      @              @      @              @      @                       @              @       @              @      �?              @      �?              @                       @      �?                      �?               @                      �?                              �?              �?                      �?      �?                      �?              �?                      @     �D@              �?     �@@              �?      4@              �?      @              �?      @                      �?              �?      @                      �?              �?      @                      @              �?                              �?                      ,@                      *@              @       @               @      @               @       @                       @               @                              @               @       @                       @               @                       @       @               @                               @              "@      &@                      @              "@      @              @      @              �?      @                      �?              �?      @              �?                              @               @                      @       @              @                               @      @      �?      @                      @      @      �?              @                              �?               @      .@     �S@       @      @      &@       @              @       @                                      @              @      @              �?      @                       @              �?      @              �?                              @              @                      $@     �P@              @      I@              @      B@              @      A@                      *@              @      5@                       @              @      3@               @       @              �?                      �?       @                       @              �?                      �?      1@              �?      .@                      "@              �?      @              �?                              @                       @              �?       @              �?                               @                      ,@              @      1@              @      �?               @                       @      �?               @                              �?               @      0@                      0@               @              @      7@      @      @      7@              @      @              @                              @                      3@                              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$�phG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�BXZ         >                  �a@�zm�4�?�           ��@       _                   �c@��֭v�?Q           0�@       ^                    @�n��)�?J            �^@       )                    �?�tU�d�?F            �]@       (                    a@E�v*��?            �J@       '                    a@a��+e�?             I@       
                     �?$��Z=;�?             F@       	                   @^@      �?              @������������������������       �                     �?������������������������       �                     �?                          �X@      �?             E@������������������������       �                     @       $                   �Z@�Kh/��?             B@                           _@     ��?             @@                           �?Z$��m�?             :@                           �?�}�+r��?
             3@������������������������       �                     &@                           \@      �?              @                          @^@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                          @_@:/����?             @������������������������       �                      @                          �]@{�G�z�?             @������������������������       �                      @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?�8��8��?             @������������������������       �                      @        !                    �?      �?             @������������������������       �                      @"       #                    �?      �?              @������������������������       �                     �?������������������������       �                     �?%       &                   @]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @*       ]                   �K@R1��HL�?'            @P@+       0                     �?��@�4Q�?&            �O@,       -                    \@�q�q�?             @������������������������       �                     �?.       /                    �?      �?              @������������������������       �                     �?������������������������       �                     �?1       R                    �?�.�?�P�?#             N@2       G                   �^@����J�?            �C@3       F                   Pb@      �?             8@4       C                    �?���y4F�?             3@5       @                   �_@*D>��?	             *@6       ?                   �^@      �?              @7       8                   `X@�8��8��?             @������������������������       �                     �?9       :                   �Y@�Q����?             @������������������������       �                      @;       <                   @[@VUUUUU�?             @������������������������       �                     �?=       >                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @A       B                    `@z�G�z�?             @������������������������       �                     @������������������������       �                     �?D       E                   p`@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @H       Q                   �d@��S���?             .@I       L                   �_@��
ц��?	             *@J       K                   �a@z�G�z�?             @������������������������       �                     @������������������������       �                     �?M       N                    ^@      �?              @������������������������       �                     @O       P                   `a@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @S       T                   `]@L�p.0�?             5@������������������������       �                     @U       \                    a@��S���?             .@V       W                   �_@���!pc�?             &@������������������������       �                     @X       [                    �?      �?             @Y       Z                   Pb@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @`       �                    �?�~�����?           �z@a       �                   Pc@�n_Y�K�?t            `h@b       q                   �i@�:v�x�?^            �c@c       d                     �?�����?             E@������������������������       �                     @e       p                   �h@��-�=��?            �C@f       g                   @_@r�q��?             8@������������������������       �                     *@h       m                   �`@���|���?             &@i       j                    b@؇���X�?             @������������������������       �                     @k       l                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?n       o                   `a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@r       u                   �Y@�͸-V<�?F            �\@s       t                    �?���Q��?             @������������������������       �                      @������������������������       �                     @v       w                   �Q@���@1�?C            �[@������������������������       �                      @x       �                    �?BMĹ��?B             [@y       ~                    `@9��8���?             8@z       {                   @]@      �?              @������������������������       �                     @|       }                   �q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?       �                   Pq@      �?             0@�       �                   `a@"pc�
�?	             &@������������������������       �                     "@������������������������       �                      @�       �                   w@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �]@Z�eY�e�?2             U@�       �                   �]@��#ۊ7�?            �C@�       �                    �?b˒�#�?            �B@�       �                   �`@�8��8��?             8@������������������������       �                     1@�       �                   �Y@����X�?             @������������������������       �                     �?�       �                   `a@r�q��?             @������������������������       �                     �?�       �                   �[@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   p@�	j*D�?             *@������������������������       �                     @������������������������       �                     "@������������������������       �                      @�       �                   �p@�����H�?            �F@�       �                    a@XB���?             =@������������������������       �        
             1@�       �                   ``@�8��8��?             (@������������������������       �                     @�       �                   �k@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                     �?      �?             0@������������������������       �                     @�       �                    a@�	j*D�?             *@�       �                   `_@      �?              @�       �                    �?z�G�z�?             @������������������������       �                     @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   t@���Q��?             @�       �                    a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   Pe@���y4F�?             C@�       �                    �?�ՙ/�?             5@�       �                   `a@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    e@��S���?	             .@������������������������       �                      @������������������������       �                     @������������������������       �        	             1@�       3                  hr@�y���?�             m@�                         0e@\��s�S�?�            �i@�       �                    �?.��Ou�?a            �c@�       �                   (r@��=�/�?,            @Q@�       �                   �`@���n(T�?+            �P@�       �                   pk@I�O���?             G@�       �                   �^@���N8�?             5@�       �                   �h@�8��8��?	             (@������������������������       �                     @�       �                   �\@z�G�z�?             @������������������������       �                     @�       �                   i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   �m@vq�-�?             9@�       �                   @]@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?���N8�?             5@�       �                    \@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �^@�<ݚ�?             2@�       �                   �a@���|���?             &@������������������������       �                     @�       �                   `c@z�G�z�?             @������������������������       �                      @�       �                   �o@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   0a@���Q��?             4@�       �                    g@r�q��?             @�       �                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?d}h���?
             ,@�       �                    �?8�Z$���?	             *@�       �                     �?"pc�
�?             &@�       �                   �a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?l��[B��?5            �U@�       �                    @�q�q�?             8@�       �                   Xp@�d�����?             3@�       �                    �?�<ݚ�?             2@�       �                   �`@      �?             0@�       �                   �]@X�<ݚ�?             "@������������������������       �                     @�       �                     �?�q�q�?             @�       �                   0m@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   l@      �?             @������������������������       �                      @�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�                          �?��~R���?&            �O@�       
                  �m@      �?             H@�                          @�q�q�?             8@�                         �l@և���X�?             5@�                           �?      �?             0@�                          �j@      �?              @������������������������       �                     �?������������������������       �                     �?                        �d@d}h���?	             ,@������������������������       �                      @                         \@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     @      	                  �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?                         @�8��8��?             8@                         a@�KM�]�?             3@                        (p@�X�<ݺ?
             2@������������������������       �                     "@                          �?�����H�?             "@                        `\@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                          �?������?	             .@������������������������       �                     @                        �_@�q�q�?             (@������������������������       �                      @                        Ph@z�G�z�?             $@������������������������       �                      @������������������������       �                      @      $                    �?�J�4�?             I@      #                  �j@�X�<ݺ?             2@                          �?      �?              @������������������������       �                     @!      "                  �i@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@%      ,                   @     ��?             @@&      '                  �e@HP�s��?             9@������������������������       �                     &@(      +                  f@؇���X�?             ,@)      *                  �]@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@-      .                   �?����X�?             @������������������������       �                     �?/      0                  @`@�q�q�?             @������������������������       �                      @1      2                  pm@      �?             @������������������������       �                      @������������������������       �                      @4      5                  �\@�����H�?             ;@������������������������       �                      @6      7                   �?`2U0*��?             9@������������������������       �                     *@8      =                   �?�8��8��?	             (@9      <                    �?r�q��?             @:      ;                  `]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @?      �                  �b@N`���}�?m             g@@      G                  �X@�9}���?Z            �c@A      F                  @h@�nkK�?             7@B      C                  @T@�C��2(�?             &@������������������������       �                     @D      E                  �U@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@H      e                  �b@>Ν�a�?M            �`@I      J                  �Y@d��z�.�?%            �N@������������������������       �                     �?K      `                  �b@��gE#�?$             N@L      M                   �?�5��	�?!            �L@������������������������       �                     *@N      O                  b@ 9�����?             F@������������������������       �                     (@P      Q                  0b@     0�?             @@������������������������       �                     @R      Y                  Po@rH��7�?             =@S      V                  `f@P���� �?             7@T      U                   �?      �?              @������������������������       �                     �?������������������������       �                     �?W      X                   @�����?             5@������������������������       �        
             3@������������������������       �                      @Z      _                   �?�8��8��?             @[      \                    �?{�G�z�?             @������������������������       �                     �?]      ^                  �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?a      b                  �b@�q�q�?             @������������������������       �                     �?c      d                   �?      �?              @������������������������       �                     �?������������������������       �                     �?f      q                  �c@h/�����?(             R@g      h                  �\@     ��?             0@������������������������       �                     @i      n                  pc@���(\��?             $@j      m                   �?z�G�z�?             @k      l                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @o      p                  ``@z�G�z�?             @������������������������       �                     �?������������������������       �                     @r      �                   �?n۶m۶�?!             L@s      |                  �_@�ӭ�a��?             B@t      u                   ]@�IєX�?             1@������������������������       �                     @v      {                  @^@�C��2(�?             &@w      z                   �?z�G�z�?             @x      y                  �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @}      �                   �?�\��N��?	             3@~                        �`@r�q��?             @������������������������       �                     �?������������������������       �                     @�      �                  `h@�	j*D�?             *@�      �                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�      �                   �?      �?             4@�      �                  �r@      �?             0@�      �                  �e@�q�q�?
             .@�      �                   _@"pc�
�?             &@������������������������       �                     @�      �                   `@���Q��?             @������������������������       �                      @������������������������       �                     @�      �                   `@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?H�$I�$�?             <@�      �                   e@"pc�
�?             &@�      �                  �c@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?�      �                   �?�IєX�?             1@�      �                  @b@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KM�KK��h[�B�&        O@     @w@     �r@     �C@     Pp@     @o@      ;@     �M@      B@      ;@     �K@      B@      @      @@      ,@      @      =@      ,@      @      =@       @              �?      �?              �?                              �?      @      <@      @              @              @      6@      @      @      6@      @      @      4@      @      �?      2@                      &@              �?      @              �?      @                      @              �?                              @               @       @      @                       @       @       @      �?               @               @              �?                      �?       @                      �?       @      @               @              �?              @                       @      �?              �?      �?                                      �?      @              �?      @                                      �?                      @              @              4@      7@      6@      4@      5@      6@      �?               @                      �?      �?              �?                      �?      �?                      3@      5@      4@      (@      *@      ,@      (@      @      @      @      @      @      @      @      �?      @      @      �?      @       @      �?              �?              @      �?      �?       @                      �?      �?      �?      �?                              �?      �?                      �?              �?                       @              @      �?              @                              �?                      �?      @              �?                              @      @                              @       @              @      @              �?      @                      @              �?                      @       @              @                      @       @                       @              @                               @      @       @      @                      @      @       @              @       @                      @              @      @              @      �?              @                              �?                       @              @                               @                      @              (@     @i@     �j@      $@     @`@     �K@      $@     �^@      9@              C@      @              @                     �A@      @              4@      @              *@                      @      @              @      �?              @                      �?      �?                      �?              �?                      �?      @                      @              �?                      .@              $@      U@      5@               @      @               @                              @      $@     �T@      2@       @                       @     �T@      2@      @      &@      "@      @      �?      @                      @      @      �?              @                              �?                      $@      @              "@       @              "@                               @              �?      @                      @              �?              @     �Q@      "@      @      ?@      @       @      ?@      @       @      6@                      1@               @      @              �?                      �?      @                      �?              �?      @                      @              �?                              "@      @                      @              "@               @                              D@      @              <@      �?              1@                      &@      �?              @                      @      �?              @                              �?              (@      @              @                      "@      @              @      �?              @      �?              @                      �?      �?              �?                              �?              @                       @      @              �?      @                      @              �?                      �?                       @      >@               @      *@              �?      @                      @              �?                      @       @                       @              @                              1@       @      R@     �c@       @     @Q@     �`@       @     �N@     @W@       @      3@      H@       @      0@      H@       @       @      B@              �?      4@              �?      &@                      @              �?      @                      @              �?      �?              �?                              �?                      "@       @      @      0@       @       @               @                               @                      @      0@              �?       @              �?                               @              @      ,@              @      @                      @              @      �?               @                       @      �?                      �?               @                              @               @      (@              @      �?               @      �?               @                              �?              @                      @      &@               @      &@               @      "@               @       @                       @               @                              @                       @              �?                      @                      E@     �F@              3@      @              ,@      @              ,@      @              (@      @              @      @              @                       @      @              �?      �?              �?                              �?              �?      @                       @              �?      �?                      �?              �?                      @                       @                              �?              @                      7@      D@              (@      B@              $@      ,@              "@      (@              @      (@              �?      �?                      �?              �?                      @      &@               @                      �?      &@              �?                              &@              @                      �?       @                       @              �?                       @      6@               @      1@              �?      1@                      "@              �?       @              �?      @              �?                              @                      @              �?                              @              &@      @              @                       @      @                       @               @       @                       @               @                       @      E@              �?      1@              �?      @                      @              �?       @                       @              �?                              $@              @      9@               @      7@                      &@               @      (@               @      @               @                              @                      "@              @       @              �?                      @       @               @                       @       @                       @               @                      @      8@               @                      �?      8@                      *@              �?      &@              �?      @              �?      @              �?                              @                      �?                      @      7@     �[@      I@      6@     @[@      9@      �?      6@              �?      $@                      @              �?      @              �?                              @                      (@              5@     �U@      9@      @     �G@      "@      �?                      @     �G@      "@      @      G@      @              *@              @     �@@      @              (@              @      5@      @                      @      @      5@      @       @      4@      �?              �?      �?              �?                              �?       @      3@                      3@               @                       @      �?      @       @      �?       @              �?               @               @       @                                       @                      �?              �?       @                      �?              �?      �?                      �?              �?              0@      D@      0@      @      @      @      @                      �?      @      @              @      �?               @      �?               @                              �?               @              �?              @      �?                                      @      "@      B@      &@      "@      :@      �?              0@      �?              @                      $@      �?              @      �?               @      �?                      �?               @                       @                      @              "@      $@              @      �?                      �?              @                      @      "@              @       @              @                               @                      @                      $@      $@              $@      @              $@      @              "@       @              @                      @       @                       @              @                      �?      @                      @              �?                              �?                      @      �?       @      9@               @      "@              �?      "@              �?                              "@              �?              �?              0@      �?              @      �?                                      @                      &@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW:+LhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�BY         �                    �?|�s;���?�           ��@       _                   �e@*`�P�?�            �w@                          `]@�aV����?N            @[@                          �_@��(\���?             D@                          �T@�8��8��?             (@                           [@��!pc�?
             &@       
                    �?�$I�$I�?             @       	                   `W@      �?             @������������������������       �                      @������������������������       �                      @                           X@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           ^@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                          �b@@4և���?             <@                           �? �q�q�?             8@                           a@�}�+r��?             3@                          �`@r�q��?             @������������������������       �                     @                          @V@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     @                          �X@      �?             @������������������������       �                     �?������������������������       �                     @       *                     �?�9���?/            @Q@        )                   �f@Y�����?             &@!       (                    b@���Q��?             $@"       #                    �?      �?              @������������������������       �                      @$       %                    Y@�q�q�?             @������������������������       �                     �?&       '                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?+       ^                   �e@&k�i}�?'             M@,       S                   �a@��hl���?%            �K@-       D                   P`@��X��?             E@.       5                   `^@@r��ճ�?             6@/       4                    I@�z�G��?             $@0       3                    �?�<ݚ�?             "@1       2                   �]@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?6       A                    �?�q�q�?             (@7       :                   �^@�<ݚ�?             "@8       9                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?;       <                   @Z@؇���X�?             @������������������������       �                     @=       >                   �_@      �?             @������������������������       �                      @?       @                    `@      �?              @������������������������       �                     �?������������������������       �                     �?B       C                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @E       R                   Pe@z�G�z�?             4@F       O                   �^@���Er�?             1@G       J                   �\@      �?             $@H       I                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @K       N                   �_@      �?             @L       M                   @E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @P       Q                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @T       U                   �b@�	j*D�?	             *@������������������������       �                     @V       W                   �]@      �?              @������������������������       �                     �?X       Y                   �c@և���X�?             @������������������������       �                      @Z       [                   Pd@z�G�z�?             @������������������������       �                     @\       ]                   pe@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @`       �                   `m@�fTx2s�?�            �p@a       t                   �i@�(>^�?@            @W@b       c                    `@4?,R��?             B@������������������������       �                     ,@d       s                   Pc@�GN�z�?             6@e       j                   0g@��s����?             5@f       g                   �[@և���X�?             @������������������������       �                     @h       i                     �?      �?             @������������������������       �                     �?������������������������       �                     @k       r                    �?@4և���?
             ,@l       q                   �`@؇���X�?             @m       n                   �\@�q�q�?             @������������������������       �                     �?o       p                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?u       |                    _@��p���?&            �L@v       {                   �a@      �?	             0@w       z                   @^@      �?              @x       y                    a@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @}       �                    `@���
8�?            �D@~       �                   �_@���Q��?             @       �                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �`@�q�q�?             B@�       �                   0a@�LQ�1	�?             7@�       �                   �Z@      �?             (@�       �                   �j@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     @�       �                   �j@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                    �?�	j*D�?
             *@�       �                    �?���Q��?             $@�       �                   0k@�q�q�?             "@������������������������       �                     @�       �                     �?���Q��?             @������������������������       �                     �?�       �                   0e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �c@��,i�?i            �e@�       �                   Pa@��?U���?Z            �b@�       �                   p@t.�eN~�?8             W@������������������������       �                     3@�       �                   �`@��L��?-            @R@�       �                   �Z@�g+�v�?             A@�       �                   `X@�g���e�?             &@�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    `@�q�q�?             "@�       �                   `q@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?�nkK�?             7@�       �                   `t@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �        	             .@�       �                   0p@�7��?            �C@������������������������       �                      @������������������������       �                    �B@�       �                   �p@<a�A���?"            �L@�       �                   @n@8��8���?             8@�       �                    b@0�����?             @�       �                   �a@r�q��?             @�       �                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    ]@�IєX�?             1@�       �                   p@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             (@�       �                   �t@�g���e�?            �@@�       �                     �?�o_��?             9@�       �                    a@�q�q�?             (@�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   @e@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?8�Z$���?             *@�       �                   �a@�q�q�?             (@������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   q@�	j*D�?             :@������������������������       �                     $@�       �                   �d@      �?	             0@������������������������       �                     @�       �                   �r@�q�q�?             (@������������������������       �                     @�       �                    f@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �c@�ل��?�            Pv@�       �                    �?(&ޏ��?             F@�       �                    \@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �? =[y��?             A@�       �                    �?      �?              @�       �                   @L@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �`@�θ�?             :@�       �                     �?���!pc�?             6@������������������������       �                      @�       �                    `@z�G�z�?             4@�       �                    `@�z�G��?             $@������������������������       �                     @�       �                    �?      �?             @�       �                   �b@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �O@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @�       �                   �\@
�ͲE�?�            �s@�       �                   �o@X�<ݚ�?             ;@�       �                    a@      �?             (@������������������������       �                     @�       �                    �?      �?              @�       �                    @:/����?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@�       2                  �j@�n�F	{�?�            �q@       	                  pf@p�h=�g�?@            @X@                          �?P���� �?             7@                        �e@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        0d@ףp=
�?             4@                         d@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             .@
                         �?���@��?1            �R@                        @g@�FVQ&�?            �@@                        �f@      �?             @������������������������       �                     �?                          �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                        @^@XB���?             =@                        i@ףp=
�?             $@                         \@      �?             @������������������������       �                     �?                        �h@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@      !                  �a@#z�i��?            �D@                        �`@��s����?             5@                        �g@      �?             0@������������������������       �                     �?������������������������       �                     .@                         @^@���Q��?             @������������������������       �                      @������������������������       �                     @"      -                  @j@      �?             4@#      $                   �?���Q��?             .@������������������������       �                     @%      (                  �f@"pc�
�?	             &@&      '                    �?      �?              @������������������������       �                     �?������������������������       �                     �?)      *                  �i@�����H�?             "@������������������������       �                     @+      ,                  @_@      �?              @������������������������       �                     �?������������������������       �                     �?.      1                   @z�G�z�?             @/      0                  �j@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @3      �                   @tA�e��?s            �g@4      Y                   �?�I	p���?g             e@5      8                  �[@JyK���?5            �U@6      7                   b@      �?             @������������������������       �                      @������������������������       �                      @9      <                  �a@U7W1�?2            �T@:      ;                  `k@�}�+r��?             3@������������������������       �                     �?������������������������       �                     2@=      B                   b@     ��?%             P@>      ?                  m@      �?              @������������������������       �                     @@      A                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @C      X                  r@4և����?!             L@D      W                   �?�4F����?            �D@E      F                  �k@^H���+�?            �B@������������������������       �                     @G      H                  �m@����e��?            �@@������������������������       �                     @I      V                  f@�q�q�?             >@J      O                  @_@����X�?             <@K      L                    �?      �?              @������������������������       �                     �?M      N                  �p@և���X�?             @������������������������       �                     @������������������������       �                     @P      U                  pd@z�G�z�?             4@Q      T                  d@������?	             .@R      S                   b@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     .@Z      �                  Xq@��SZ�$�?2            @T@[      �                   b@�vp��?$            �J@\      e                  �]@l&{��?!            �H@]      b                   �?      �?	             (@^      a                  �[@z�G�z�?             @_      `                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @c      d                  `\@����X�?             @������������������������       �                     @������������������������       �                      @f      w                  �`@����>�?            �B@g      r                  q@7�ٔ_�?             =@h      k                  pk@      �?             8@i      j                  �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?l      q                  pb@���N8�?             5@m      n                  �_@�����H�?             "@������������������������       �                     @o      p                  0m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@s      t                    �?���Q��?             @������������������������       �                     �?u      v                   �?      �?             @������������������������       �                     @������������������������       �                     �?x                         �?      �?              @y      z                   �?����X�?             @������������������������       �                     �?{      |                  Pa@�q�q�?             @������������������������       �                     �?}      ~                  �d@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                  `]@      �?             <@������������������������       �                     @�      �                    �?�q�q�?             8@�      �                  8r@��.k���?             1@������������������������       �                      @������������������������       �                     "@�      �                   �?����X�?             @�      �                  �a@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                    �?؇���X�?             5@������������������������       �                      @�      �                   �?�}�+r��?
             3@�      �                  �o@      �?              @������������������������       �                     @�      �                  �q@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�t�b�      h�h(h+K ��h-��R�(KM�KK��h[�B(&        F@     �w@     �s@      B@     @n@     �X@      6@      K@     �@@      @      @@      @      @      @       @      @      @       @      @       @      �?       @       @                       @               @                       @              �?                      �?       @                              @      �?              @                              �?              �?                      :@       @              7@      �?              2@      �?              @      �?              @                      �?      �?                      �?              �?                      *@                      @                      @      �?                      �?              @              2@      6@      =@      @      �?      @      @              @      @              @                       @      @               @      �?                      @               @                       @      @                       @                              �?              (@      5@      9@      "@      5@      9@      "@      (@      5@      @      &@      @              @      @               @      @               @      @               @                              @                      �?              �?              @       @               @      @              �?      �?              �?                              �?              �?      @                      @              �?      @                       @              �?      �?              �?                              �?               @      �?                      �?               @                      @      �?      ,@      @      �?      &@      @              @       @              @       @                                      @      @              �?      �?              �?      �?                                      �?       @                              �?      @              �?                              @                      @              "@      @              @                      @      @                      �?              @      @                       @              @      �?              @                      �?      �?                      �?              �?              @                      ,@     �g@     �P@      @     �M@      ?@              ?@      @              ,@                      1@      @              1@      @              @      @              @                      �?      @              �?                              @              *@      �?              @      �?               @      �?              �?                      �?      �?              �?                              �?              @                      @                              �?      @      <@      :@               @      ,@               @      @              �?      @                      @              �?                      �?                               @      @      :@      (@      @       @               @      �?               @                              �?              �?      �?              �?                              �?                      8@      (@              4@      @              "@      @              �?       @              �?                               @               @      �?              @                      @      �?                      �?              @                      &@                      @      "@              @      @              @      @                      @              @       @                      �?              @      �?              @                              �?              �?                              @      &@      `@     �A@      &@     @^@      1@      "@     @T@       @              3@              "@      O@       @      @      9@       @      @      @      �?      �?              �?                      �?      �?                      @      @               @      @                      @               @                      @                              6@      �?              @      �?              @                              �?              .@               @     �B@               @                             �B@               @      D@      .@      �?      5@       @      �?      @      �?              @      �?              @      �?              @                              �?              �?              �?                              0@      �?              @      �?              @                              �?              (@              �?      3@      *@      �?      &@      *@              @      @               @      @               @                              @              @      �?              @                              �?      �?      @       @              @       @                       @              @              �?                               @                       @      2@                      $@               @       @                      @               @      @              @                       @      @                      @               @               @     �`@     �j@      �?      <@      .@              �?      "@              �?                              "@      �?      ;@      @      �?      @              �?      @                      @              �?                              �?                      4@      @              0@      @                       @              0@      @              @      @              @                      @      @              @       @                       @              @                              �?              "@      �?              "@                              �?              @              @     �Z@      i@      @      2@      @      @      @      @                      @      @      @       @      @       @       @               @       @                       @               @              @                              �?                      .@              @      V@     @h@      �?      2@     �S@      �?       @      4@      �?               @      �?                                       @               @      2@               @      @               @                              @                      .@              0@      M@               @      ?@              �?      @                      �?              �?       @                       @              �?                      �?      <@              �?      "@              �?      @                      �?              �?       @                       @              �?                              @                      3@              ,@      ;@              @      1@              �?      .@              �?                              .@              @       @                       @              @                      $@      $@              @      "@              @                       @      "@              �?      �?              �?                              �?              �?       @                      @              �?      �?              �?                              �?              @      �?               @      �?                      �?               @                       @              @     �Q@      ]@      @      J@     @\@              7@      P@               @       @               @                               @              5@      O@              �?      2@              �?                              2@              4@      F@              @      �?              @                       @      �?                      �?               @                      *@     �E@              *@      <@              *@      8@                      @              *@      4@              @                      $@      4@               @      4@              @      @              �?                      @      @                      @              @                      @      0@              @      &@               @      &@                      &@               @                       @                              @               @                              @                      .@      @      =@     �H@      @      .@     �A@      @      (@      A@              @      @              @      �?              �?      �?                      �?              �?                      @                       @      @                      @               @              @      @      <@      @      @      7@              @      5@               @      �?               @                              �?              �?      4@              �?       @                      @              �?       @              �?                               @                      (@      @               @                      �?      @              �?      @                                      �?              @      @               @      @                      �?               @      @              �?                      �?      @              �?                              @              �?                      @      �?                      �?              @                      ,@      ,@              @                      $@      ,@               @      "@               @                              "@               @      @              �?      @              �?                              @              �?                      2@      @                       @              2@      �?              @      �?              @                      @      �?                      �?              @                      &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF<KdhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�Bc         �                  �c@�p"��?�           ��@       �                   u@0%̘��?�           Ȅ@       �                   �`@4yۓǉ�?�           ��@       �                    �?ġ�]+��?�            `p@       Z                    �?�M=-\�?�            �h@       Y                   �t@Ɯ��2��?^            �a@       N                   �p@F3r����?]            `a@                            �?,"dM�?M            �]@	                           �?X�Cc�?             ,@
                          �`@�	j*D�?             *@                          0k@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?       -                   `_@4�b$���?F            @Z@                          `X@p=
ףp�?             D@������������������������       �                      @       *                   �_@(������?             C@                           �?�n#،A�?             A@                          0i@ףp=
�?             $@                          `g@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @       )                   �^@      �?             8@       "                   `\@��uJ���?             3@       !                   �^@.y0��k�?             *@                           �?�8��8��?             (@������������������������       �                     @                            [@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?#       (                    I@VUUUUU�?             @$       %                    �?      �?             @������������������������       �                     �?&       '                   `]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @+       ,                    `@      �?             @������������������������       �                     @������������������������       �                     �?.       /                   �`@`��>�b�?,            @P@������������������������       �                     5@0       9                   @a@4_�g���?             F@1       8                    �?և���X�?             @2       7                   �m@      �?             @3       6                    W@      �?             @4       5                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?:       M                   �p@b˒�#�?            �B@;       <                    �?,R�n��?             B@������������������������       �                     @=       J                   @c@     ��?             @@>       C                   �a@ĳ���o�?             >@?       @                    ^@�θ�?             *@������������������������       �                     "@A       B                   Pl@      �?             @������������������������       �                     @������������������������       �                     �?D       E                   �^@�IєX�?
             1@������������������������       �                     *@F       I                    �?      �?             @G       H                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @K       L                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?O       P                   q@��Q��?             4@������������������������       �                     @Q       X                    \@������?             1@R       W                   c@X�<ݚ�?             "@S       V                    Z@����X�?             @T       U                   hr@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                      @[       �                    �?�S����?%            �L@\       i                     �?�������?             F@]       b                   @_@�.�?��?
             .@^       _                    �?�����H�?             "@������������������������       �                     @`       a                   `i@�q�q�?             @������������������������       �                      @������������������������       �                     �?c       f                    @      �?             @d       e                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?g       h                   �p@      �?             @������������������������       �                     �?������������������������       �                     @j       o                   @[@�%d���?             =@k       n                   �k@����X�?             @l       m                    W@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @p       {                   �_@ˠT�x�?             6@q       r                   �Z@�m۶m��?
             ,@������������������������       �                     �?s       z                   `^@8�Z$���?	             *@t       u                    �?����X�?             @������������������������       �                     �?v       w                    �?r�q��?             @������������������������       �                      @x       y                   n@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @|       }                   �\@      �?              @������������������������       �                     @~       �                   0d@���Q��?             @       �                   `@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @�	j*D�?             *@�       �                    �?"pc�
�?             &@�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �W@؇���X�?             @������������������������       �                     @�       �                     �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    _@     @�?*             P@�       �                    �?޾�z�<�?             *@�       �                    \@�����H�?             "@������������������������       �                     @�       �                     �?r�q��?             @������������������������       �                     �?�       �                    �?z�G�z�?             @�       �                    X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   `]@      �?             @������������������������       �                      @������������������������       �                      @�       �                   0j@8��(y��?"            �I@�       �                   �^@�_[��?             ?@�       �                   @^@0�����?             5@�       �                   �h@     @�?             0@�       �                   `]@/����?             ,@�       �                   @b@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                   �a@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   �a@�z�G��?             $@�       �                   `@���Q��?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     4@�       �                    �?�E�4���?�            �w@�       �                    �?     q�?M             `@�       �                   Pc@�Ö�jw�?=            �X@�       �                   �l@ƇG+���?&            �O@�       �                   �k@���|���?            �@@�       �                    �?y0��k��?             :@�       �                   a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �]@�8��8��?             8@������������������������       �                     @�       �                   �a@�ՙ/�?             5@�       �                   h@������?             1@������������������������       �                     (@�       �                    �?z�G�z�?             @�       �                   �j@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   `g@      �?             @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    ]@j�Y�H��?             >@�       �                    �?      �?              @������������������������       �                      @�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?�0�~�4�?             6@�       �                   0b@�X�<ݺ?             2@������������������������       �        
             0@�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    a@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?����X�?            �A@�       �                    p@:ɨ��?            �@@������������������������       �        	             *@�       �                   �r@      �?             4@�       �                   �d@      �?             (@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   0f@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    f@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   0m@ףp=
��?             >@�       �                    Y@Z�K8�?             :@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �j@��+��?             5@�       �                   @W@~h����?
             ,@�       �                   �`@Y�����?             &@�       �                     �?      �?              @������������������������       �                      @�       �                   �d@      �?             @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       "                   �?`{�>α�?�             o@�                          �?�~����?            �E@�                           �?A�F<��?             C@                         �`@      �?             (@                        `o@����X�?             @������������������������       �                      @������������������������       �                     @                         b@���Q��?             @                        `a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @	                         �?y0��k��?             :@
                        �p@      �?              @������������������������       �                     @                        �r@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         @�)O�?             2@                        �`@     ��?
             0@                        p@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?                        j@���Q��?             @������������������������       �                     �?                         b@      �?             @                        �n@�q�q�?             @������������������������       �                     �?                        �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @      !                   @z�G�z�?             @                         �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @#      F                    �?��+$�?|            �i@$      A                  �e@�-���?#             I@%      6                  �`@��P���?            �D@&      -                  �c@\-��p�?             =@'      (                  �_@      �?             0@������������������������       �                     "@)      ,                   n@؇���X�?             @*      +                  �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @.      /                  �i@�θ�?             *@������������������������       �                     @0      1                  �c@�z�G��?             $@������������������������       �                      @2      3                  �d@      �?              @������������������������       �                     @4      5                  �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @7      @                  �d@�q�q�?	             (@8      ?                   @      �?              @9      :                  0a@      �?             @������������������������       �                      @;      >                  �a@      �?             @<      =                  p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @B      E                  �e@X�<ݚ�?             "@C      D                   �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @G      H                  �G@���B���?Y            �c@������������������������       �                     @I      p                  �b@@�0�!��?X             c@J      g                   �?V��z4�?'             O@K      f                   �?�q�q�?             H@L      a                   @8����?             G@M      N                  Pa@�G�z�?             D@������������������������       �                     .@O      `                   b@�q�����?             9@P      U                  �g@և���X�?             5@Q      R                  �a@r�q��?             @������������������������       �                     @S      T                   �?      �?              @������������������������       �                     �?������������������������       �                     �?V      ]                   �?������?             .@W      X                  �a@z�G�z�?             $@������������������������       �                     �?Y      \                  b@�����H�?             "@Z      [                  �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @^      _                  `b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @b      c                  @`@r�q��?             @������������������������       �                     @d      e                  �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @h      i                   `@d}h���?	             ,@������������������������       �                     @j      k                  p`@�z�G��?             $@������������������������       �                      @l      o                   �?      �?              @m      n                  pb@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @q      �                   @|)����?1            �V@r      u                  �O@(�s���?-             U@s      t                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?v      �                   �?H�!b	�?+            @T@w      �                  pd@ >�֕�?%            �Q@x      �                  Pd@<���D�?            �@@y      �                   q@`Jj��?             ?@z      �                   �?ףp=
�?             4@{      �                  Hp@�KM�]�?
             3@|                         c@�X�<ݺ?	             2@}      ~                  �\@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                      @������������������������       �                    �B@������������������������       �                     &@�      �                   �?և���X�?             @�      �                  �f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�      �                  �\@���B���?             :@�      �                   \@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                  �]@؇���X�?             5@������������������������       �                     @�      �                   �?r�q��?	             2@�      �                  @_@�θ�?             *@������������������������       �                     �?�      �                   �?r�q��?             (@�      �                    �?�C��2(�?             &@������������������������       �                     @�      �                  0`@      �?             @������������������������       �                      @�      �                  v@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?��?���?0            @Q@�      �                  h@�z�G��?             D@�      �                    �?�z�G��?             $@�      �                  �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?����X�?             @������������������������       �                      @�      �                   V@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                    �?��S���?             >@�      �                   �?      �?              @�      �                   c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                   f@8�A�0��?             6@�      �                  �^@�t����?             1@�      �                  pl@�C��2(�?             &@�      �                  �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�      �                  �d@�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                  �q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                   �?�%d���?             =@�      �                  @^@0�����?             2@������������������������       �                     @�      �                   g@��!pc�?             &@�      �                  �_@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KM�KK��h[�Bx*        C@     `v@      u@      A@     `s@     t@      A@     r@     �s@      7@     �e@     �P@      3@     �`@     �G@      1@     �Z@      2@      1@     �Z@      0@      $@     @W@      0@              "@      @              "@      @              @      @              @                              @              @                              �?      $@      U@      &@       @      <@      @       @                      @      <@      @      @      ;@      @              "@      �?              @      �?              @                              �?              @              @      2@      @      @      *@      @      �?      &@      �?      �?      &@                      @              �?      @              �?                              @                              �?       @       @       @       @               @                      �?       @              �?       @                                      �?               @                      @              @      �?              @                              �?               @      L@      @              5@               @     �A@      @              @      @              @      @              �?      @              �?      �?                      �?              �?                               @               @                      �?               @      ?@      @       @      ?@      @              @               @      ;@      @      �?      :@      @              $@      @              "@                      �?      @                      @              �?              �?      0@                      *@              �?      @              �?      �?              �?                              �?                       @              �?      �?                      �?              �?                                      �?      @      *@              @                      @      *@              @      @               @      @               @      �?               @                              �?                      @               @                               @                               @       @      :@      =@       @      1@      9@      �?      @      "@              �?       @                      @              �?       @                       @              �?              �?      @      �?              �?      �?              �?                              �?      �?      @              �?                              @              �?      (@      0@              @       @               @       @               @                               @              @              �?      @      ,@      �?       @      &@      �?                               @      &@               @      @              �?                      �?      @                       @              �?      @                      @              �?                              @              @      @              @                       @      @               @      �?               @                              �?                       @              "@      @              "@       @              @      �?              @                              �?              @      �?              @                      @      �?                      �?              @                               @      @      D@      4@      �?       @      $@      �?               @                      @      �?              @                      �?      �?              @      �?              �?                      �?      �?                                      @               @       @                       @               @              @      C@      $@      @      2@      $@      @      .@      @      @      $@      @      �?      $@      @              "@      �?              "@                              �?      �?      �?       @      �?      �?              �?                              �?                               @       @                              @                      @      @              @       @              �?       @                       @              �?                       @                              @              4@              &@     @]@      o@      @      K@     �P@       @     �E@     �J@       @     �@@      <@      �?      $@      6@      �?      $@      .@              �?      �?              �?                              �?      �?      "@      ,@              @              �?      @      ,@              @      *@                      (@              @      �?              @      �?                      �?              @                      �?              �?       @      �?      �?              �?      �?                                      �?               @                              @      �?      7@      @              @      @                       @              @       @                       @              @              �?      3@       @      �?      1@                      0@              �?      �?              �?                              �?                       @       @                       @               @                      $@      9@              $@      7@                      *@              $@      $@              "@      @              �?       @              �?                               @               @      �?               @                              �?              �?      @                      @              �?                               @      @      &@      ,@      @      @      ,@      @              �?      @                                      �?      �?      @      *@      �?      @      @      �?      @      @      �?      �?      @                       @      �?      �?      @      �?      �?              �?                              �?                              @              @                      @                              @              @              @     �O@     �f@      @      4@      3@      @      4@      .@       @      @      @               @      @               @                              @       @      @               @      �?                      �?               @                               @              �?      .@      $@              �?      @                      @              �?       @              �?                               @      �?      ,@      @      �?      (@      @      �?      $@                      $@              �?                               @      @              �?                      �?      @              �?       @                      �?              �?      �?              �?                              �?                      �?               @              �?              @      �?              �?      �?                                      �?                      @             �E@     `d@              *@     �B@              "@      @@              @      9@              �?      .@                      "@              �?      @              �?       @                       @              �?                              @              @      $@                      @              @      @               @                      �?      @                      @              �?       @              �?                               @              @      @              @      @              @      @                       @              @      �?              �?      �?                      �?              �?                       @                       @                              @              @      @              @       @                       @              @                              @              >@     �_@              @                      ;@     �_@              3@     �E@              0@      @@              ,@      @@              *@      ;@                      .@              *@      (@              "@      (@              @      �?              @                      �?      �?                      �?              �?                      @      &@               @       @              �?                      �?       @              �?       @                       @              �?                              @               @      @                      @               @                      @                      �?      @                      @              �?       @                       @              �?                       @                      @      &@                      @              @      @               @                      �?      @              �?       @              �?                               @                      @               @     �T@              @     �S@              �?       @                       @              �?                      @     @S@              @     �P@              @      =@               @      =@               @      2@               @      1@              �?      1@              �?      @                      @              �?                              *@              �?                              �?                      &@               @                             �B@                      &@              @      @              �?      @                      @              �?                       @                      5@      @              @       @              @                               @              2@      @              @                      .@      @              $@      @                      �?              $@       @              $@      �?              @                      @      �?               @                      �?      �?              �?                              �?                      �?              @              @      H@      1@      @      5@      0@      @      @              �?       @              �?                               @               @      @                       @               @      @                      @               @                              ,@      0@              �?      @              �?      @              �?                              @                      @              *@      "@              (@      @              $@      �?              �?      �?              �?                              �?              "@                       @      @                      @               @                      �?      @                      @              �?              �?      ;@      �?      �?      0@      �?              @              �?      "@      �?              "@      �?                      �?              "@              �?                              &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJؽ�hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�d         �                   P`@R�
\��?�           ��@       �                    �?������?�            u@                             �?�4���?�            @o@                          r@~K紂�?            �I@                           _@     ��?             @@                           Z@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@	                          �k@�$�_�?             3@
                          ``@r�q��?             (@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@                          `[@؇���X�?             @������������������������       �                     @                           b@      �?             @������������������������       �                     �?                          �^@�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                           ]@�d�����?	             3@������������������������       �                      @                           �?@�0�!��?             1@������������������������       �                      @                           �?�q�q�?             "@                          @e@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @!       j                    _@pHZ���?x            �h@"       #                    Q@����ۊ�?a             d@������������������������       �                     �?$       W                    �?      �?`             d@%       &                    [@�v��"��?C            �\@������������������������       �                     @'       R                   @]@T��2�7�?A            �[@(       O                   �\@��n&��?-            @T@)       6                    �?�j���?*            @S@*       +                   �g@hE#߼�?
             .@������������������������       �                     @,       3                   �a@�g���e�?             &@-       2                    �?      �?              @.       1                   �^@      �?             @/       0                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @4       5                   q@�q�q�?             @������������������������       �                      @������������������������       �                     �?7       L                    s@"����?              O@8       E                   �`@����0L�?            �M@9       :                   �X@4��hZ�?             =@������������������������       �                     *@;       <                   @Y@     ��?             0@������������������������       �                     @=       D                   �[@$�q-�?	             *@>       C                   �_@r�q��?             @?       @                   �Z@�q�q�?             @������������������������       �                     �?A       B                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @F       K                   @U@(;L]n�?             >@G       H                   �S@r�q��?             @������������������������       �                     @I       J                    c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@M       N                   �t@�q�q�?             @������������������������       �                     �?������������������������       �                      @P       Q                    �?      �?             @������������������������       �                      @������������������������       �                      @S       T                   @g@(;L]n�?             >@������������������������       �        	             .@U       V                   j@��S�ۿ?             .@������������������������       �                     �?������������������������       �        
             ,@X       Y                   �^@��'����?             G@������������������������       �                      @Z       c                   �b@0�/5mv�?             C@[       b                   �`@h�����?             <@\       ]                   �_@      �?              @������������������������       �                     @^       _                    �?z�G�z�?             @������������������������       �                     @`       a                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@d       i                   �q@      �?             $@e       h                    S@r�q��?             @f       g                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @k       x                    �?�S����?             C@l       s                   0`@�m۶m��?             <@m       r                    �?������?	             .@n       q                   `_@d}h���?             ,@o       p                   �a@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?t       u                   0a@8�Z$���?             *@������������������������       �                     "@v       w                    k@      �?             @������������������������       �                      @������������������������       �                      @y       z                    �?�Q����?             $@������������������������       �                      @{       |                   �_@      �?              @������������������������       �                      @}       ~                   P`@�q�q�?             @������������������������       �                      @       �                    `@      �?             @������������������������       �                      @������������������������       �                      @�       �                   @d@T|d�O_�?;            �U@�       �                   �[@z�c��?5            �R@�       �                    �?L]n���?             >@������������������������       �                     �?�       �                     �?П[;U��?             =@������������������������       �                     �?�       �                   `R@H�$I�$�?             <@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �Z@T���N@�?             9@������������������������       �                     .@�       �                    �?��(\���?             $@�       �                    [@      �?              @������������������������       �                     �?�       �                   �\@؇���X�?             @������������������������       �                     @�       �                   �K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �_@�2(&��?!             F@�       �                    s@�Cc}h��?             <@�       �                    �?      �?             8@�       �                   �k@     @�?             0@�       �                    �?�n���?             "@�       �                     �?      �?              @������������������������       �                     �?�       �                   @c@:/����?             @�       �                   @Y@�8��8��?             @�       �                   `]@      �?             @������������������������       �                     �?�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                     �?؇���X�?             @������������������������       �                     �?�       �                   @p@r�q��?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?             @�       �                   �|@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                     �?      �?	             0@������������������������       �                      @�       �                   `c@և���X�?             ,@�       �                   �a@�n_Y�K�?             *@�       �                    `@�eP*L��?             &@�       �                   @_@և���X�?             @�       �                   �[@���Q��?             @������������������������       �                     �?������������������������       �      �?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@�       �                   @E@z����?�            �x@�       �                    �?h3�݃��?            �A@�       �                    Y@��|���?             6@�       �                   �G@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �`@�IєX�?             1@������������������������       �                     �?�       �                   �a@     ��?             0@������������������������       �                     @�       �                     �?H�z�G�?	             $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   pc@      �?              @�       �                   Pb@      �?             @������������������������       �                     �?�       �                   `]@VUUUUU�?             @������������������������       �                     �?�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   b@��
ц��?             *@�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @�       �                     @�q�q�?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �?����G�?�            �v@�       S                  �b@�'�W
�?�            Pt@�       N                  �c@p=
ףp�?X            �a@�       M                   c@��4`��?T            �`@�                          �?�}�X���?S            ``@�                         hp@���%�3�?&             O@�                         Hp@mdk����?             E@�       �                   pf@�^�����?            �C@�       �                   �a@{�G�z�?             @�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @�                         `n@�M���?             A@�       �                     �?"	��p�?             =@������������������������       �                     �?�                         �m@/�����?             <@�                         �a@5���?             :@�                         �k@��JÝ�?             7@�                         `a@������?             1@�                          �`@�q�q�?             @�       �                   @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                        �a@؇���X�?             ,@������������������������       �                     @                         ]@      �?              @                         [@      �?              @������������������������       �                     �?������������������������       �                     �?      	                  @_@r�q��?             @������������������������       �                     @
                         �?      �?              @������������������������       �                     �?������������������������       �                     �?                        Pl@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @                         �?P���Q�?             4@������������������������       �        
             3@������������������������       �                     �?      >                  pa@ٜSu��?-            @Q@      =                   �?H.�!���?              I@                          �?�%^�?            �E@                         �?��S�ۿ?             .@                        �\@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@      $                   �?X�Cc�?             <@       !                  l@      �?             @������������������������       �                     �?"      #                  �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @%      4                  �_@�q�q�?             8@&      +                  �a@��
ц��?
             *@'      (                   �?z�G�z�?             @������������������������       �                      @)      *                  Pi@�q�q�?             @������������������������       �                      @������������������������       �                     �?,      -                  �j@      �?              @������������������������       �                     @.      3                   _@      �?             @/      0                  0b@�q�q�?             @������������������������       �                     �?1      2                  0m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?5      6                  �a@"pc�
�?             &@������������������������       �                     @7      8                   �?���Q��?             @������������������������       �                      @9      <                  �`@�q�q�?             @:      ;                  �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @?      J                  @b@D�n�3�?             3@@      A                  `a@      �?             0@������������������������       �                     @B      I                    �?�q�q�?             "@C      H                  �r@և���X�?             @D      E                  �k@z�G�z�?             @������������������������       �                      @F      G                  p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @K      L                  �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @O      P                  `a@�8��8��?             @������������������������       �                      @Q      R                  �e@      �?             @������������������������       �                     @������������������������       �                     �?T      w                   �?BBF����?t             g@U      \                  `\@X�Cc�?#             L@V      W                  �Z@z�G�z�?             .@������������������������       �                     �?X      Y                  �[@؇���X�?             ,@������������������������       �                     @Z      [                   o@      �?              @������������������������       �                      @������������������������       �                     @]      h                    �?v�2t5�?            �D@^      _                  `c@���|���?	             &@������������������������       �                     �?`      g                  �e@�z�G��?             $@a      b                  `]@�<ݚ�?             "@������������������������       �                     �?c      f                  `o@      �?              @d      e                  @n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?i      v                  �f@*;L]n�?             >@j      k                  `k@8�A�0��?             6@������������������������       �                     @l      u                   d@     ��?
             0@m      n                  �d@X�Cc�?             ,@������������������������       �                     @o      p                  Pe@      �?              @������������������������       �                     @q      r                  �_@���Q��?             @������������������������       �                      @s      t                  ``@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @x      y                  �c@�e$´�?Q             `@������������������������       �                     �?z      �                  �p@     P�?P             `@{      �                  �c@|<SvL�?7             W@|      �                  �l@�-^~Z�?4            @V@}      �                  �\@���U�?             �L@~                        �h@؇���X�?             @������������������������       �                     �?������������������������       �                     @�      �                  i@p���?             I@�      �                  `^@���7�?             6@�      �                  �c@r�q��?             @������������������������       �                     @�      �                   g@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@������������������������       �                     <@�      �                  d@      �?             @@������������������������       �                     .@�      �                  �d@V��6���?             1@�      �                  Pd@      �?             @�      �                    �?�q�q�?             @������������������������       �                     �?�      �                  �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                  @e@8�Z$���?
             *@�      �                  �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �f@ףp=
�?             $@������������������������       �                     @�      �                  �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                  �f@tk~X��?             B@�      �                  @r@��hJ,�?             A@�      �                  �d@      �?             $@�      �                   �?�q�q�?             @������������������������       �                      @�      �                   �?      �?             @������������������������       �                      @������������������������       �                      @�      �                  @`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     8@������������������������       �                      @�      �                    �?t����{�?            �B@�      �                  @q@؇���X�?             @������������������������       �                     @�      �                  �s@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  0f@.�?�P��?             >@�      �                  �f@3������?             =@������������������������       �                     @�      �                  �h@9��8���?             8@������������������������       �                     @�      �                   a@��[r��?             5@�      �                  0l@�.�?��?             .@�      �                   a@�$I�$I�?             @������������������������       �                      @�      �                  �_@{�G�z�?             @������������������������       �                      @�      �                  Pi@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �^@      �?              @�      �                  0m@�q�q�?             @������������������������       �                     �?�      �                  �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?r�q��?             @�      �                  �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�t�b�P     h�h(h+K ��h-��R�(KM�KK��h[�B8+        F@     0w@     �s@      <@     �m@      R@      (@      f@     �N@      �?      7@      ;@      �?      "@      6@              �?      (@              �?                              (@      �?       @      $@               @      $@               @      �?               @                              �?                      "@      �?      @                      @              �?      @                      �?              �?       @              �?      �?                      �?              �?                              �?                      ,@      @                       @              ,@      @               @                      @      @               @      @                      @               @                      @              &@     @c@      A@      @     @`@      :@                      �?      @     @`@      9@      @     �X@      (@                      @      @     �X@      "@      @     @Q@       @      @     �P@      @      �?      &@      @              @              �?      @      @      �?      @      �?      �?      @      �?      �?              �?                      �?      �?                              @                       @                      �?       @                       @              �?              @      L@      @       @      K@      @      �?      9@      @              *@              �?      (@      @                      @      �?      (@              �?      @              �?       @                      �?              �?      �?              �?                              �?                      @                      @              �?      =@              �?      @                      @              �?      �?                      �?              �?                              8@              �?       @              �?                               @                       @       @               @                               @              =@      �?              .@                      ,@      �?                      �?              ,@              �?      @@      *@                       @      �?      @@      @      �?      ;@              �?      @                      @              �?      @                      @              �?      �?                      �?              �?                              4@                      @      @              �?      @              �?       @                       @              �?                              @              @              @      8@       @      @      6@       @      @      &@              @      &@              @      @                      @              @                              @              �?                              &@       @              "@                       @       @                       @               @               @       @      @                       @       @       @      @               @               @              @                       @       @               @       @                                       @      0@      N@      &@      0@     �G@      &@      @      9@       @      �?                       @      9@       @                      �?       @      9@      �?      �?       @              �?                               @              �?      7@      �?              .@              �?       @      �?      �?      @      �?      �?                              @      �?              @                      @      �?                      �?              @                       @              *@      6@      "@      @      ,@      "@      @      (@      "@       @      @      "@       @      @      @       @      @      @                      �?       @      @       @      �?      @       @      �?      �?       @      �?                              �?       @                       @              �?                       @              �?                              �?                      �?      @                      �?              �?      @                      @              �?       @              �?                               @      �?      @              �?                              @               @       @               @      �?               @                              �?                      �?               @       @                       @               @      @               @      @              @      @              @      @              @       @              �?                       @       @                       @              @      �?                      �?              @                       @                              �?                      *@              0@     �`@     �n@      @      3@      &@      @      *@      @      @      �?                      �?              @                      �?      (@      @                      �?      �?      (@      @              @              �?      @      @              �?      �?              �?                              �?      �?      @       @      �?      �?       @                      �?      �?      �?      �?                      �?      �?      �?              �?                              �?                      @                      @      @               @      @                      @               @                      @       @              �?       @                       @              �?                      @              &@     �\@     �m@      "@      X@     �k@      @     �O@     �Q@      @      O@      Q@      @      O@     @P@      @     �E@      .@      @      8@      ,@      @      8@      &@       @      �?       @              �?      �?              �?                              �?       @              �?                      �?       @                       @      7@      "@       @      2@      "@              �?               @      1@      "@       @      1@      @       @      1@      @              *@      @              �?       @              �?      �?                      �?              �?                              �?              (@       @              @                      @       @              �?      �?              �?                              �?              @      �?              @                      �?      �?                      �?              �?               @      @               @                              @                              @                       @              @                              @              3@      �?              3@                              �?              3@      I@              &@     �C@              &@      @@              �?      ,@              �?      @                      @              �?                              &@              $@      2@               @       @                      �?               @      �?                      �?               @                       @      0@              @      @              @      �?               @                       @      �?               @                              �?               @      @                      @               @       @              �?       @                      �?              �?      �?                      �?              �?                      �?                       @      "@                      @               @      @                       @               @      �?              �?      �?                      �?              �?                      �?                              @               @      &@              @      $@                      @              @      @              @      @              @      �?               @                       @      �?                      �?               @                               @               @                       @      �?                      �?               @                              @      @      �?       @                       @      @      �?              @                              �?               @     �@@     �b@              4@      B@              @      (@              �?                       @      (@                      @               @      @               @                              @              1@      8@              @      @              �?                      @      @               @      @              �?                      �?      @              �?       @                       @              �?                              @              �?                      *@      1@              *@      "@              @                      @      "@              @      "@                      @              @      @              @                       @      @                       @               @      �?               @                              �?               @                               @       @      *@     �\@              �?               @      (@     �\@       @      @     @U@       @      @     �T@               @     �K@              �?      @              �?                              @              �?     �H@              �?      5@              �?      @                      @              �?       @                       @              �?                              0@                      <@       @       @      <@                      .@       @       @      *@               @       @              �?       @                      �?              �?      �?              �?                              �?              �?               @              &@      �?               @      �?                                       @      �?              "@                      @      �?               @      �?                                       @              �?       @                       @              �?                      @      =@              @      =@              @      @               @      @                       @               @       @               @                               @              @      �?              @                              �?                      8@               @               @      3@      0@              @      �?              @                       @      �?                      �?               @               @      *@      .@       @      *@      ,@                      @       @      *@      "@              @               @      $@      "@      �?      @      "@      �?      @       @               @              �?       @       @               @              �?               @      �?                                       @              �?      @              �?       @                      �?              �?      �?              �?                              �?                      @      �?      @              �?       @                       @              �?                              @                              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJX��vhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�^         �                   p`@��j�`�?�           ��@       o                    i@�i15v�?�             t@       F                    �?@{}^�D�?f            �c@       A                   �_@�mc���?@            @Y@                           `@������?<            �W@                          @^@��=��*�?            �B@                           �?t=9%�R�?             ;@       	                     �?�(\����?
             4@������������������������       �                     �?
                          @Z@�lO���?	             3@                          �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@                          `]@�$I�$I�?             @                          �S@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �Z@      �?             @������������������������       �                     �?������������������������       �                     @                           �?p=
ףp�?             $@                           [@�$I�$I�?             @                          �_@      �?             @                          `Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @       0                   b@P*�n���?'             M@        #                   �Y@�����H�?             B@!       "                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @$       %                   �`@`Jj��?             ?@������������������������       �        
             1@&       '                     �?؇���X�?
             ,@������������������������       �                     �?(       /                    �?8�Z$���?	             *@)       .                   �T@�8��8��?             (@*       -                    a@      �?              @+       ,                   `]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?1       @                    �?"pc�
�?             6@2       3                     �?�S����?             3@������������������������       �                      @4       7                   @U@�IєX�?             1@5       6                   �S@�q�q�?             @������������������������       �                     �?������������������������       �                      @8       ;                    �?�m۶m��?	             ,@9       :                    _@      �?              @������������������������       �                     @������������������������       �                      @<       ?                   c@r�q��?             @=       >                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @B       C                   0`@�8��8��?             @������������������������       �                     @D       E                   �X@�q�q�?             @������������������������       �                      @������������������������       �                     �?G       R                   `[@�X�C�?&             L@H       Q                   `c@B{	�%��?             2@I       N                    �?�"�O�|�?             1@J       M                    \@�����H�?             "@K       L                   @Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @O       P                   `]@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?S       d                   `_@&:~�Q�?             C@T       ]                    _@Y�����?             6@U       \                    ^@      �?             (@V       W                   �Y@      �?              @������������������������       �                     @X       Y                    \@      �?             @������������������������       �                      @Z       [                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @^       a                   �_@ףp=
��?             $@_       `                   �Z@r�q��?             @������������������������       �                     �?������������������������       �                     @b       c                   �[@      �?             @������������������������       �                     �?������������������������       ��q�q�?             @e       l                    �?     ��?             0@f       g                    ^@����X�?
             ,@������������������������       �                     @h       k                   �N@      �?              @i       j                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @m       n                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?p       �                    �?�,�-v(�?j            �d@q       ~                    Z@�xRvQ��?K            @]@r       u                   �W@��1+��?             ;@s       t                   �x@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?v       y                    �?b�r���?	             .@w       x                   @]@�q�q�?             @������������������������       �                      @������������������������       �                     @z       }                   �n@�q�q�?             "@{       |                   �X@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       �                   �k@���S�Y�?:            �V@�       �                   @Z@�(�I�8�?             =@������������������������       �                      @�       �                   �\@PN��T'�?             ;@�       �                    �?�X�<ݺ?	             2@������������������������       �                     0@�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?             "@������������������������       �                     @�       �                     �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   pb@�h�*��?+            �N@�       �                   �\@�(\����?             D@�       �                   �Z@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �A@�       �                   �o@:/����?             5@������������������������       �                     &@�       �                   �d@�Q����?             $@�       �                   `c@{�G�z�?             @�       �                    �?VUUUUU�?             @�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    \@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �`@�q�q��?             H@�       �                    �?�����?             3@�       �                    �?�E��ӭ�?             2@�       �                    �?r�q��?             @�       �                   Xp@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   @r@�q�q�?             (@�       �                     �?�����H�?             "@�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    g@��Θ���?             =@�       �                    _@ܶm۶m�?             <@�       �                    �?�nkK�?             7@�       �                   @\@�8��8��?             (@������������������������       �                     @�       �                   �\@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�                          �?(Ll�٧�?           �y@�                         Pc@�M��?_            �c@�       �                   0m@��#[���?@            �Y@�       �                    �?BݪxF�?"            �I@�       �                   �k@:/����?             E@�       �                   �k@0\�Uo��?             C@�       �                    �?��aE�?            �A@�       �                    �?Q�a�r��?             >@�       �                   �a@���(\��?             $@�       �                   �Y@����X�?             @������������������������       �                     �?�       �                   �i@r�q��?             @������������������������       �                     @�       �                   @j@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �g@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @_@R���Q�?             4@�       �                   �]@{�G�z�?             $@�       �                   �W@�8��8��?             @������������������������       �                     �?�       �                   �a@���Q��?             @������������������������       �                     �?�       �                   Pb@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   Pa@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    b@�z�G��?             $@�       �                   �e@�<ݚ�?             "@�       �                    U@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   `b@���Q��?             @������������������������       �                     �?�       �                   �b@      �?             @������������������������       �                     �?�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �e@�<ݚ�?             "@�       �                   pb@���Q��?             @�       �                   `b@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    ]@�Ƽ����?            �I@�       �                   �b@      �?             ,@�       �                   �r@�z�G��?             $@�       �                    �?      �?             @�       �                   �n@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �q@@0.1�r�?            �B@������������������������       �                     5@�                          �r@     ��?	             0@������������������������       �                     �?                        �a@�r����?             .@                        `a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     &@                        `T@H �6��?            �K@      
                   �?      �?              @      	                  �e@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                          �?TnH/h]�?            �G@                         �?     ��?             0@                        `a@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @                         _@��a�n`�?             ?@                         �?      �?             $@                        �p@X�<ݚ�?             "@                         �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                        �i@�����?             5@                        �c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        
             1@      �                   �?��S%���?�            �o@       K                   �?RSv���?�            `k@!      F                   �?t����?@            �Z@"      5                  c@�r����?6            �V@#      *                  �^@¦	^_�?             ?@$      '                    �?      �?             (@%      &                  �n@և���X�?             @������������������������       �                     @������������������������       �                     @(      )                  �f@���Q��?             @������������������������       �                      @������������������������       �                     @+      2                  �q@�S����?             3@,      -                   �?      �?             0@������������������������       �                     �?.      1                    �?��S�ۿ?
             .@/      0                  @b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@3      4                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @6      E                  �`@����˵�?$            �M@7      <                   �?��<D�m�?            �H@8      9                  �d@      �?              @������������������������       �                     �?:      ;                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @=      >                    �?��Y��]�?            �D@������������������������       �                     0@?      D                  @^@`2U0*��?             9@@      C                  �j@�}�+r��?
             3@A      B                   g@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@������������������������       �                     @������������������������       �                     $@G      H                    �?      �?
             0@������������������������       �                     $@I      J                  �k@r�q��?             @������������������������       �                     @������������������������       �                     �?L      S                  �a@�}��_�?I            @\@M      N                   �?���7�?             6@������������������������       �                     0@O      R                  p`@r�q��?             @P      Q                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @T      a                  �b@p�-@�Z�?:            �V@U      X                   �?"pc�
�?
             6@V      W                  �o@z�G�z�?             @������������������������       �                     @������������������������       �                     �?Y      Z                  �b@@�0�!��?             1@������������������������       �                     @[      \                  @e@�z�G��?             $@������������������������       �                     @]      `                  @_@      �?             @^      _                  0m@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?b      �                  e@�?�0���?0            @Q@c      d                  �[@z�5���?             C@������������������������       �                     @e      f                  `]@,\&p��?             ?@������������������������       �                     @g      �                  �d@pƵHPS�?             :@h      s                  �c@�8��8��?             8@i      l                    �?h/�����?             "@j      k                  �b@      �?              @������������������������       �                     �?������������������������       �                     �?m      r                  `a@������?             @n      o                  �p@�Q����?             @������������������������       �                     @p      q                  �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @t      {                   �?hE#߼�?             .@u      v                   g@�8��8��?             @������������������������       �                     �?w      z                  8r@���Q��?             @x      y                  pd@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @|      }                    �?�����H�?             "@������������������������       �                      @~                         a@؇���X�?             @������������������������       �                     @�      �                  �i@�q�q�?             @������������������������       �                     �?�      �                  d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                  �s@�n`���?             ?@�      �                   f@r�q��?             >@�      �                  �e@�d�����?             3@�      �                  �j@@�0�!��?             1@�      �                  0g@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     (@������������������������       �                      @������������������������       �                     &@������������������������       �                     �?�      �                  �^@�Kh/���?             B@������������������������       �                     @�      �                    �?�v�`��?             ?@�      �                   �?�q�q�?             @������������������������       �                     �?�      �                  �c@z�G�z�?             @������������������������       �                      @�      �                  @q@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   a@���H�?             9@������������������������       �                     �?�      �                  �p@r�q��?             8@�      �                  Pa@�M�]��?             1@������������������������       �                      @�      �                  �c@���ĳ��?             .@�      �                   �?z�G�z�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                  `d@���Q��?             $@�      �                  d@r�q��?             @�      �                  �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                  �`@      �?             @�      �                  �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B�(       �P@     �v@     �r@     �F@      k@      N@      @@      W@     �@@      1@     @P@      3@      ,@      P@      1@      $@      4@      @      @      3@      @       @      1@      �?              �?               @      0@      �?       @              �?                      �?       @                              0@              �?       @      @               @      �?               @                              �?      �?              @      �?                                      @      @      �?       @      @      �?       @      �?      �?       @      �?      �?              �?                              �?                               @      @                      @                      @      F@      $@              @@      @              @       @                       @              @                      =@       @              1@                      (@       @              �?                      &@       @              &@      �?              @      �?               @      �?               @                              �?              @                      @                              �?      @      (@      @      @      (@      @                       @      @      (@      �?       @      �?                      �?               @                       @      &@      �?       @      @                      @               @                              @      �?               @      �?               @                              �?              @                              @      @      �?       @      @                              �?       @                       @              �?              .@      ;@      ,@       @      ,@       @      �?      ,@       @      �?       @              �?       @                       @              �?                              @                      @       @                       @              @              �?                      *@      *@      (@      (@       @       @      "@              @      @              @      @                      �?              @                       @      �?              �?      �?                                      �?      @                      @       @      @              �?      @              �?                              @      @      �?              �?                       @      �?              �?      &@      @              $@      @              @                      @      @               @      @               @                              @               @              �?      �?              �?                              �?              *@     @_@      ;@      (@      X@      "@      @      1@      @      �?      &@                      &@              �?                      @      @      @      @               @                       @      @                              @      @              �?      @              �?                              @              @              @     �S@      @      @      7@       @                       @      @      7@              �?      1@                      0@              �?      �?                      �?              �?                      @      @                      @              @       @                       @              @                      @      L@       @      �?     �C@              �?      @              �?                              @                     �A@               @      1@       @              &@               @      @       @       @      �?       @      �?      �?      �?              �?      �?                      �?              �?              �?                      �?              �?      �?                                      �?              @              �?      =@      2@              @      *@              @      *@              �?      @              �?       @              �?                               @                      @              @       @              �?       @              �?      �?              �?                              �?                      @              @                      �?              �?      7@      @      �?      7@      @      �?      6@              �?      &@                      @              �?      @              �?                              @                      &@                      �?      @                      @              �?                              �?      5@     �b@     `n@      2@     @S@      O@      &@      P@      ;@      $@      7@      2@      $@      0@      0@      $@      0@      (@      @      0@      (@      @      *@      (@      �?      @      @               @      @              �?                      �?      @                      @              �?       @              �?                               @      �?       @              �?                               @              @      "@      @      @       @      @      �?       @      @      �?                               @      @              �?                      �?      @                      @              �?              @              �?                      �?      @                              @      @              @       @               @       @               @                               @              @                              �?       @      @              �?                      �?      @                      �?              �?       @              �?                               @              @                                      @              @       @              @       @              @      �?                      �?              @                              �?              @              �?     �D@      "@              @      @              @      @              @      @              �?      @              �?                              @               @                      @                              @      �?      A@       @              5@              �?      *@       @      �?                              *@       @               @       @               @                               @              &@              @      *@     �A@       @      @               @      @                      @               @                              @              @      @     �A@      @              &@      @              @                      @      @                                      @              @      8@              @      @              @      @              �?      @                      @              �?                      @                              �?               @      3@               @       @               @                               @                      1@      @     �Q@     �f@       @      J@     �d@              *@     @W@              (@     �S@              "@      6@              @      @              @      @                      @              @                      @       @                       @              @                      @      0@              �?      .@                      �?              �?      ,@              �?       @              �?                               @                      (@               @      �?                      �?               @                      @      L@              @      G@               @      @              �?                      �?      @              �?                              @              �?      D@                      0@              �?      8@              �?      2@              �?       @                       @              �?                              0@                      @                      $@              �?      .@                      $@              �?      @                      @              �?               @     �C@      R@              �?      5@                      0@              �?      @              �?       @                       @              �?                              @       @      C@     �I@              2@      @              @      �?              @                              �?              ,@      @              @                      @      @              @                      @      @              @       @                       @              @                              �?       @      4@     �G@       @      ,@      6@                      @       @      ,@      .@              @               @      "@      .@       @      @      .@      �?      @      @              �?      �?                      �?              �?              �?      @      @      �?      �?      @                      @      �?      �?              �?                              �?                       @              �?      @      &@      �?       @      @      �?                               @      @               @      �?               @                              �?                       @              �?       @                       @              �?      @                      @              �?       @                      �?              �?      �?                      �?              �?                       @                      @      9@              @      9@              @      ,@              @      ,@              @       @                       @              @                              (@               @                              &@              �?              �?      3@      0@                      @      �?      3@      &@              @       @                      �?              @      �?               @                       @      �?               @                              �?      �?      .@      "@                      �?      �?      .@       @      �?       @       @               @              �?      @       @      �?              @      �?              �?                      �?      �?                                      @              @      @              @      �?               @      �?               @                              �?              @                      �?      @              �?      �?              �?                              �?                       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���EhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�BXa         d                   �?�:���?�           ��@       �                    �?z,�p���?x           X�@       �                   �c@6f�1��?�            `s@                            �?�n�z���?�            �p@                          @_@��s����?             E@                          @b@      �?             (@       
                    �?�q�q�?             "@       	                   �`@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @                           f@��S�ۿ?             >@                           �?`2U0*��?             9@������������������������       �                     $@                          �`@��S�ۿ?
             .@                          @Z@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@                          �g@z�G�z�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       K                   pg@�X�c�?�             l@       @                   P`@�6��O�?/            �T@                          �Z@� �)��?$            �M@������������������������       �                     @       5                    �?|��?���?#             K@       4                   �d@ k U��?            �A@        3                   �f@     `�?             @@!       "                   @R@N�s�-�?             ?@������������������������       �                      @#       .                   `_@4��hZ�?             =@$       '                    �?p=
ףp�?             $@%       &                   �T@      �?             @������������������������       �                     �?������������������������       �                     @(       -                    I@      �?             @)       *                   @[@      �?             @������������������������       �                     �?+       ,                    ]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @/       0                    �?�}�+r��?             3@������������������������       �                     �?1       2                   @e@�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?������������������������       �                     �?������������������������       �                     @6       7                    `@R��Xp�?
             3@������������������������       �                     @8       ?                   0d@������?             .@9       >                   �b@���Q��?             $@:       ;                   �]@؇���X�?             @������������������������       �                     @<       =                   pa@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @A       B                    Y@t���?             7@������������������������       �                     �?C       D                    �?��2(&�?
             6@������������������������       �                     �?E       J                    �?�����?	             5@F       G                   pf@�r����?             .@������������������������       �                     $@H       I                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @L       M                   �X@¥@7�g�?[            �a@������������������������       �                     �?N       �                   0c@���3`��?Z            �a@O       p                   �l@�K���8�?P            �_@P       S                   �Y@:/����?#             L@Q       R                   �j@      �?             @������������������������       �                     �?������������������������       �                     @T       g                    �?޾�z�<�?              J@U       \                   �j@z��V�k�?            �E@V       W                   �[@���N8�?             5@������������������������       �                      @X       Y                    `@�n_Y�K�?             *@������������������������       �                     @Z       [                   0b@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @]       b                   �_@��2(&�?             6@^       _                   �k@�q�q�?             @������������������������       �                     @`       a                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?c       f                   @\@      �?	             0@d       e                   �[@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @h       o                   0l@x�5?,�?             "@i       l                   �j@      �?              @j       k                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?m       n                    `@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?q       z                    �?�����?-            �Q@r       y                   @^@8߄*�u�?             1@s       t                   Pn@0�����?             @������������������������       �                     @u       v                   �Z@      �?             @������������������������       �                      @w       x                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@{       |                   �]@��B�<�?             �J@������������������������       �                     ,@}       �                    �?���	7I�?            �C@~       �                   @_@�B��j��?            �@@       �                   �`@      �?              @������������������������       �                     @�       �                   �p@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �`@`2U0*��?             9@�       �                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     4@�       �                   �_@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?���Q��?
             .@������������������������       �                     �?�       �                   �[@/����?	             ,@������������������������       �                     @�       �                   Pd@      �?              @������������������������       �                      @�       �                   �^@      �?             @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    g@      �?             @�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    s@����!p�?             F@�       �                   Pe@vKQ#�?            �A@�       �                   a@p=
ףp�?             4@�       �                   (p@X�Cc�?             ,@�       �                   Pi@      �?             $@������������������������       �                      @�       �                   @`@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   `o@      �?             @������������������������       �                     @�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     �?�r����?
             .@������������������������       �                     �?�       �                   �r@؇���X�?	             ,@������������������������       �                     (@������������������������       �                      @������������������������       �                     "@�       G                  �d@r<��+��?�            Pq@�       �                    �?�������?�            �i@�       �                     �?�G�z��?6             T@�       �                   �`@����X�?             5@������������������������       �        	             &@�       �                   �a@���Q��?             $@�       �                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   `X@rfg�Ka�?&            �M@������������������������       �                     @�       �                   `_@n۶m۶�?$             L@�       �                    �?� �	��?             9@������������������������       �                     @�       �                    d@b�2�tk�?             2@�       �                    �?��S���?             .@�       �                   �h@      �?             ,@�       �                   �[@      �?             @������������������������       �                     �?�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �a@���Q��?             $@������������������������       �                      @�       �                   �l@      �?              @������������������������       �                     @�       �                   �\@�q�q�?             @������������������������       �                     �?�       �                   �o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   @_@tH�����?             ?@�       �                   �b@      �?             @�       �                   �]@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @b@`2U0*��?             9@������������������������       �                     2@�       �                    c@؇���X�?             @�       �                   `q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �_@H��M��?T             _@�       �                   �\@R��Xp�?             3@������������������������       �                     @�       �                    �?{�G�z�?             .@�       �                   �`@���(\��?             $@�       �                   @L@z�G�z�?             @�       �                   `P@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     @�       �                   @]@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @���Q��?             @�       �                   P`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �Y@VR�s&�?F            @Z@������������������������       �                     @�       2                   a@H��'�?C            @Y@�       +                   @P��!�?.            @R@�       *                  �d@     8�?'             P@�                           �?�Z&rA��?%             M@�                         �q@�d�����?             3@�                         �n@     ��?
             0@�       �                    _@�q�q�?             "@������������������������       �                     �?�                          �a@      �?              @������������������������       �                     @                         �?���Q��?             @                        c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @      
                   �?�q�q�?             @      	                  `]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?      )                  �c@<KQ�^��?            �C@                         �?��)�8�?             A@                         \@H�z�G�?             $@������������������������       �                      @                        �^@      �?              @������������������������       �                     @                        `o@      �?              @������������������������       �                     �?������������������������       �                     �?                        �]@�q�q�?             8@������������������������       �                     @                        `@�G��l��?             5@������������������������       �                     @                         j@b�2�tk�?             2@                        `^@�<ݚ�?             "@������������������������       �                     �?                        d@      �?              @������������������������       �                     �?������������������������       �                     @      $                  @_@X�<ݚ�?             "@       !                  �l@���Q��?             @������������������������       �                      @"      #                  0m@�q�q�?             @������������������������       �                      @������������������������       �                     �?%      &                  `a@      �?             @������������������������       �                     �?'      (                  l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @,      -                  �`@�<ݚ�?             "@������������������������       �                     @.      1                  �i@�q�q�?             @/      0                  �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @3      @                  Pl@�S�r
^�?             <@4      7                  @^@      �?	             (@5      6                  pk@�q�q�?             @������������������������       �                     @������������������������       �                      @8      9                  @f@�8��8��?             @������������������������       �                     �?:      ?                   �?���Q��?             @;      <                  `a@      �?             @������������������������       �                     �?=      >                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?A      B                  �p@      �?             0@������������������������       �                     "@C      F                    �?և���X�?             @D      E                  @t@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @H      S                   �?�nr���?1            @R@I      R                  0f@d}h���?             ,@J      K                  @^@�q�q�?             "@������������������������       �                     @L      Q                    �?���Q��?             @M      N                   �?      �?             @������������������������       �                      @O      P                  Pe@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @T      a                  @g@=H��?&            �M@U      `                  @^@��2����?#            �K@V      ]                  pl@�;�;�?             :@W      \                    �?��S�ۿ?             .@X      Y                  �i@      �?              @������������������������       �                     @Z      [                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @^      _                  Pe@���!pc�?             &@������������������������       �                     @������������������������       �                      @������������������������       �                     =@b      c                  Pn@      �?             @������������������������       �                      @������������������������       �                      @e      �                  �c@Ɉ�F�(�?X            `b@f      �                  �c@`�ĪW��?F             ]@g      |                  `]@ �`�B�?>            �Y@h      {                   �?K&:~��?             3@i      p                  �Y@     @�?             0@j      k                    �?�q�q�?             @������������������������       �                     �?l      o                   �?z�G�z�?             @m      n                  `X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @q      r                  �Z@���(\��?             $@������������������������       �                     �?s      z                   �?x�5?,�?             "@t      w                   \@      �?              @u      v                  �]@      �?              @������������������������       �                     �?������������������������       �                     �?x      y                   Y@�q�q�?             @������������������������       �                      @������������������������       �      �?             @������������������������       �                     �?������������������������       �                     @}      �                   �?,��3S��?2            �T@~      �                   �?�8��8��?             H@      �                  �_@VR�s&�?            �A@�      �                  �]@�G�z�?             4@�      �                   �?����X�?             @�      �                  q@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  �b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                  @a@8�Z$���?             *@�      �                   b@r�q��?             (@�      �                   ^@�C��2(�?             &@�      �                  �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�      �                  `r@�r����?	             .@������������������������       �                     (@�      �                   u@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?/y0��k�?	             *@������������������������       �                     @�      �                  @V@z�G�z�?             $@������������������������       �                      @������������������������       �                      @�      �                   c@Z��;҂�?            �A@�      �                   `@     0�?             @@�      �                  �a@:/����?             5@������������������������       �                     (@�      �                  �i@h/�����?             "@�      �                   Y@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �                   �?��!pc�?             &@�      �                  xr@x�5?,�?             "@�      �                  �`@      �?              @������������������������       �                     @�      �                  `a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                  �e@@4և���?             ,@�      �                    �?      �?              @�      �                  �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                  @d@`Jj��?             ?@�      �                  �[@�t����?             1@������������������������       �                     "@�      �                  `]@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     ,@�t�b��     h�h(h+K ��h-��R�(KM�KK��h[�B�)       �L@      w@     0s@      B@     �q@     �p@      6@     �h@     @V@      5@     `g@      M@              A@       @              @      @              @      @              @      @              @                              @                      @              @                      <@       @              8@      �?              $@                      ,@      �?              @      �?                      �?              @                      "@                      @      �?              �?      �?                      �?              �?                      @              5@      c@      I@      &@     �C@      @@      $@      B@      *@                      @      $@      B@       @      @      9@      @      @      9@      @      @      9@      @                       @      @      9@      �?       @      @      �?      �?      @              �?                              @              �?      @      �?      �?       @      �?      �?                               @      �?               @                              �?               @              �?      2@                      �?              �?      1@                      1@              �?                                      �?      @                      @      &@      @      @                              &@      @              @      @              @      �?              @                      �?      �?                      �?              �?                              @              @              �?      @      3@      �?                              @      3@              �?                       @      3@               @      *@                      $@               @      @                      @               @                              @      $@     �\@      2@                      �?      $@     �\@      1@      @      Z@      0@      @     �D@      &@              �?      @              �?                              @      @      D@       @      @     �A@      @              0@      @               @                       @      @              @                      @      @                      @              @              @      3@               @      @                      @               @      �?               @                              �?              �?      .@              �?      @                      @              �?                               @              �?      @      @      �?      @       @              �?       @                       @              �?              �?      @              �?                              @                              �?       @     �O@      @      �?      .@      �?      �?      @      �?              @              �?       @      �?               @              �?              �?      �?                                      �?              $@              �?      H@      @              ,@              �?      A@      @      �?      =@      @              @      @              @                      �?      @              �?                              @      �?      8@              �?      @                      @              �?                              4@                      @      �?              @                              �?      @      $@      �?      �?                      @      $@      �?              @              @      @      �?       @                      �?      @      �?              �?      �?                      �?              �?              �?      @              �?      �?              �?                              �?                       @              �?      (@      ?@      �?      (@      6@      �?      $@      "@              "@      @              @      @               @                      @      @                      @              @                      @              �?      �?      @                      @      �?      �?              �?                              �?                       @      *@                      �?               @      (@                      (@               @                              "@      ,@     �U@      f@      "@     �T@     @\@      �?      9@      K@              @      .@                      &@              @      @               @      @               @                              @              @              �?      3@     �C@              @              �?      0@     �C@              ,@      &@              @                      @      &@              @       @              @      @              �?      @                      �?              �?       @              �?                               @              @      @                       @              @       @              @                      �?       @                      �?              �?      �?                      �?              �?                              �?                      @      �?       @      <@      �?      �?      @      �?              @                      @      �?                              �?      �?              �?                              �?              �?      8@                      2@              �?      @              �?       @                       @              �?                              @       @     �L@     �M@      @      &@      @              @              @      @      @      @      @      �?      @      �?              @      �?                      �?              @                      �?                              @      �?              @                      �?      �?                      �?              �?                       @      @              �?      @                      @              �?                      �?              @      G@     �K@                      @      @      G@     �I@      �?      ?@     �D@      �?      8@     �C@      �?      2@     �C@              @      ,@              @      *@              @      @              �?                       @      @                      @               @      @               @      �?               @                              �?                       @                      @               @      �?              �?      �?              �?                              �?              �?              �?      *@      9@      �?      *@      4@      �?      @      @               @              �?      �?      @                      @      �?      �?                      �?              �?                              $@      ,@                      @              $@      &@              @                      @      &@               @      @              �?                      �?      @              �?                              @              @      @              @       @               @                      �?       @                       @              �?                       @       @                      �?               @      �?               @                              �?                      @              @                      @       @              @                      @       @              �?       @              �?                               @              @              @      .@      $@      @      @      @       @              @                      @       @                      �?      @       @      �?                              @       @               @       @                      �?               @      �?               @                              �?              �?                      (@      @              "@                      @      @              @      �?              @                              �?                      @      @      @      P@              @      &@              @      @                      @              @       @              @      �?               @                      �?      �?              �?                              �?                      �?                      @      @      �?     �J@      @      �?     �I@      @      �?      6@              �?      ,@              �?      @                      @              �?       @              �?                               @                      @      @               @      @                                       @                      =@       @               @                       @       @                      5@     @U@     �D@      5@      L@     �C@      5@     �K@      :@      "@      "@      �?      @      "@      �?       @      @              �?                      �?      @              �?       @                       @              �?                               @              @      @      �?      �?                      @      @      �?      @      @              �?      �?              �?                              �?               @      @                       @               @       @                              �?      @                      (@      G@      9@      @      6@      5@       @      4@      *@       @      @      &@       @      @              �?      �?                      �?              �?                      �?      @                      @              �?                               @      &@               @      $@              �?      $@              �?      @                      @              �?                              @              �?                              �?              *@       @              (@                      �?       @                       @              �?              @       @       @      @                               @       @               @                               @      @      8@      @      @      5@      @       @      1@       @              (@               @      @       @       @               @                       @       @                              @              @      @       @      @      @      �?      @       @      �?      @                               @      �?                      �?               @                      �?                      �?      �?                      �?              �?                      @                      �?      *@              �?      @              �?      �?                      �?              �?                              @                      @              =@       @              .@       @              "@                      @       @                       @              @                      ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:9)bhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�B�e         �                  ht@�;NWR�?�           ��@       5                  c@9�m13�?�           ��@       �                   `_@(D(hV�?5            @       m                    �?S[S���?l            �d@       <                   `@h/�����?Z             b@       5                   @^@jM��?/            �R@       
                     �?     ��?(             P@       	                   @\@z�G�z�?             @������������������������       �                     �?������������������������       �                     @       "                    \@$ΕCQ��?#            �M@                          �Z@Έ����?             9@                           �?�q-��?             *@������������������������       �                     @                          `X@ףp=
��?             $@������������������������       �                     �?                          �Y@�n���?             "@                           �?:/����?             @                           �?���Q��?             @������������������������       �                     �?                          �\@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @                           \@      �?              @������������������������       �                     �?������������������������       �                     �?       !                    ]@�q�q�?             (@                           �?      �?              @������������������������       �                      @                            �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @#       0                    �?�g+�v�?             A@$       -                    �?8����?             7@%       ,                   �_@�����?             3@&       +                    �?������?
             1@'       *                   pj@z�G�z�?             @(       )                   @\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                      @.       /                    Y@      �?             @������������������������       �                      @������������������������       �      �?              @1       2                    k@"pc�
�?             &@������������������������       �                      @3       4                   �W@�q�q�?             @������������������������       �                      @������������������������       �                     �?6       ;                    �?Y�����?             &@7       8                    �?�$I�$I�?             @������������������������       �                     �?9       :                   �\@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @=       V                    �?�?�� ��?+            @Q@>       E                   @Y@z5�h$�?             >@?       D                   @E@      �?             @@       A                    Y@�q�q�?             @������������������������       �                     �?B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?F       U                   �n@R�}e�.�?             :@G       T                   `m@�q�q�?             8@H       S                   �k@�E��ӭ�?             2@I       N                   `i@     ��?
             0@J       K                   �\@�C��2(�?             &@������������������������       �                     @L       M                   pf@z�G�z�?             @������������������������       �                     �?������������������������       �                     @O       R                   �\@���Q��?             @P       Q                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @W       j                   �b@�e����?            �C@X       c                   0m@�'�`d�?            �@@Y       b                   b@�����H�?             2@Z       [                   �g@�<ݚ�?             "@������������������������       �                     �?\       ]                   Pk@      �?              @������������������������       �                     @^       _                     �?z�G�z�?             @������������������������       �                     @`       a                   `a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@d       e                   �\@�q�q�?
             .@������������������������       �                     @f       g                   0n@r�q��?             (@������������������������       �                     �?h       i                   `b@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?k       l                   Po@      �?             @������������������������       �                     @������������������������       �                     @n                           �?�p�F�:�?             7@o       ~                    �?&%�ݒ��?             5@p       y                   �`@.k��\�?             1@q       r                   `]@.y0��k�?
             *@������������������������       �                     @s       t                    X@0�����?             @������������������������       �                     @u       v                     �?VUUUUU�?             @������������������������       �                     �?w       x                    �?      �?              @������������������������       �                     �?������������������������       �                     �?z       }                   �]@      �?             @{       |                   `X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��*e���?�            �t@�       �                   �a@�g\��?"             J@�       �                   q@HP�s��?             9@������������������������       �                     7@������������������������       �                      @�       �                    �?@�����?             ;@�       �                   �`@�ӭ�a��?             2@�       �                   p@$�q-�?	             *@������������������������       �                      @�       �                   `b@z�G�z�?             @������������������������       �                      @�       �                   q@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   Ph@���Q��?             @������������������������       �                     �?�       �                   �a@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   `@X�<ݚ�?             "@������������������������       �                     @�       �                   Pb@z�G�z�?             @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   0`@�ܴND��?�            pq@�       �                     �?�Np���?k            �d@�       �                    �?�X�C�?	             ,@�       �                     @��8��8�?             (@�       �                    �?�q�q�?             "@�       �                   @l@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   `n@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   0j@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   @s@K����?b             c@�       �                   q@0\K5���?^            �b@�       �                    f@���{�?T            �`@�       �                   �a@�2����?R            @`@�       �                   �p@*񎴠��?/            �Q@�       �                    �?��eP*L�?.            �P@�       �                   �O@Ļ��|�?              G@�       �                   `R@z�G�z�?             4@������������������������       �                     �?�       �                    �?�S����?             3@�       �                    [@      �?             (@�       �                   �_@և���X�?             @������������������������       �                      @�       �                   �`@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    `@�K8��?             :@�       �                    \@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�x?r���?             6@�       �                   0k@�E�_���?             5@�       �                   �`@r�q��?             @������������������������       �                      @�       �                   �a@      �?             @�       �                   k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?��S�ۿ?	             .@�       �                   �`@�C��2(�?             &@������������������������       �                     @�       �                   0l@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   �k@�G�z��?             4@�       �                    @��8��8�?	             (@�       �                    �?p=
ףp�?             $@�       �                    �?�$I�$I�?             @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�G�z�?#             N@�       �                   �i@�����?             E@�       �                   Pd@�q�q�?             (@�       �                   @^@z�G�z�?             $@������������������������       �                     @�       �                   `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     >@�       �                    �?�)O�?             2@�       �                   `j@      �?              @�       �                   @\@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     @������������������������       �        
             ,@�       �                   @]@���Q��?             @������������������������       �                     @������������������������       �                      @�                          �? �Cc��?<             \@�                         0g@FSӂU��?            �H@�                         �`@�d�����?
             3@                         �`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                         U@@4և���?             ,@������������������������       �                      @                        �e@r�q��?             @������������������������       �                     �?������������������������       �                     @                        �a@ĳ���o�?             >@	      
                  �p@���7�?             6@������������������������       �                     .@                          �?؇���X�?             @������������������������       �                     @                        Pa@      �?             @������������������������       �                     @������������������������       �                     �?                         a@      �?              @������������������������       �                     �?                        �b@0�����?             @                         �?      �?             @                        k@      �?              @������������������������       �                     �?������������������������       �                     �?                        �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @      "                    �?��~R���?            �O@                         �?X�Cc�?             ,@                         a@�q�q�?             @������������������������       �                     @������������������������       �                      @       !                  �r@      �?              @������������������������       �                     @������������������������       �                     �?#      0                  b@����X�?            �H@$      -                   �?�חF�P�?             ?@%      *                   �?�<ݚ�?	             2@&      )                  �`@d}h���?             ,@'      (                  �h@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @+      ,                  �a@      �?             @������������������������       �                     @������������������������       �                     �?.      /                  Xr@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?1      2                  @e@      �?             2@������������������������       �                     @3      4                  �b@�	j*D�?             *@������������������������       �                     @������������������������       �                     "@6      �                   @�L�B���?~            �g@7      F                  �O@j�V��?w             f@8      A                  �e@&�q-�?
             *@9      :                   �?�q�q�?             "@������������������������       �                      @;      <                   ^@և���X�?             @������������������������       �                      @=      @                   �?z�G�z�?             @>      ?                  �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @B      C                   �?      �?             @������������������������       �                      @D      E                  �[@      �?              @������������������������       �                     �?������������������������       �                     �?G      �                   �?�av��?m            `d@H      a                   �?nb��G|�?d            �b@I      \                  `e@R���Q�?             D@J      Y                  �d@�i�V��?             6@K      P                  pc@     ��?             0@L      M                  �p@���Q��?             @������������������������       �                      @N      O                  �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?Q      V                  d@��!pc�?             &@R      S                  hp@�����H�?             "@������������������������       �                     @T      U                  �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?W      X                   n@      �?              @������������������������       �                     �?������������������������       �                     �?Z      [                  �r@r�q��?             @������������������������       �                     @������������������������       �                     �?]      `                  Pm@�X�<ݺ?             2@^      _                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@b      �                  @g@�;��t��?J            @[@c      �                  `@&��`�?H            �Z@d      u                    �?fN~K$e�?#             G@e      l                   �?�t����?             1@f      k                   �?�C��2(�?             &@g      h                  �d@�q�q�?             @������������������������       �                     �?i      j                  �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @m      t                  �p@�q�q�?             @n      o                  �\@z�G�z�?             @������������������������       �                     �?p      s                  @^@      �?             @q      r                   k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?v      }                  �[@4�����?             =@w      x                  @[@և���X�?             @������������������������       �                      @y      z                  �m@z�G�z�?             @������������������������       �                     @{      |                  �q@      �?              @������������������������       �                     �?������������������������       �                     �?~      �                  �n@8�A�0��?             6@      �                  �^@ףp=
��?             $@�      �                   �?      �?              @������������������������       �                     �?�      �                   �?և���X�?             @�      �                  �m@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�      �                  `]@r�q��?	             (@�      �                  `\@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?�����H�?             "@�      �                  `e@      �?              @�      �                  �d@      �?             @������������������������       �                      @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   �?P���Q�?%             N@�      �                    �? ���J��?            �C@�      �                  �q@z�G�z�?             @�      �                  �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     A@�      �                    �?�����?             5@�      �                  �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �l@�X�<ݺ?
             2@������������������������       �                     *@�      �                  Pd@z�G�z�?             @������������������������       �                      @�      �                  `e@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  �i@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             ,@�      �                   �?և���X�?             ,@�      �                   d@r�q��?             @������������������������       �                     �?������������������������       �                     @�      �                  �c@      �?              @������������������������       �                     @������������������������       �                     @�      �                   �?v[X���?             G@�      �                   �?���k���?            �@@�      �                  v@8�Z$���?             :@������������������������       �                     $@�      �                   �?      �?             0@������������������������       �                     @�      �                  �]@���Q��?             $@������������������������       �                     @�      �                    �?և���X�?             @������������������������       �                      @�      �                  @b@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                  ``@؇���X�?             @������������������������       �                     @�      �                   �?�q�q�?             @�      �                   y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                   u@�	j*D�?             *@������������������������       �                     �?�      �                  �]@      �?             (@������������������������       �                     @�      �                  pc@և���X�?             @������������������������       �                      @�      �                  @|@z�G�z�?             @�      �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KM�KK��h[�B�+        L@     Pw@     s@     �K@      u@     �r@      H@     �r@     @c@      <@     �Q@      Q@      :@      Q@      I@      5@     �C@      .@      1@      C@      "@              �?      @              �?                              @      1@     �B@      @      $@      (@      @      @      @      @      @                       @      @      @              �?               @      @      @       @      @       @       @      @                      �?               @       @                       @               @                                       @              �?      �?                      �?              �?              @      @              @      @                       @              @      �?                      �?              @                              @              @      9@       @      @      0@              @      *@              @      *@              @      �?              �?      �?              �?                              �?              @                              (@               @                      �?      @                       @              �?      �?                      "@       @               @                      �?       @                       @              �?              @      �?      @      @      �?       @              �?              @               @      @                                       @                      @      @      =@     �A@       @      3@      "@       @               @       @              �?      �?                      �?              �?                      �?      �?                                      �?              3@      @              3@      @              *@      @              *@      @              $@      �?              @                      @      �?                      �?              @                      @       @              �?       @              �?                               @               @                               @              @                               @      @      $@      :@              @      :@               @      0@               @      @              �?                      �?      @                      @              �?      @                      @              �?      �?                      �?              �?                              "@              @      $@              @                       @      $@              �?                      �?      $@                      $@              �?              @      @                      @              @                       @      @      2@      �?      @      1@      �?      @      *@      �?      �?      &@                      @      �?      �?      @                      @      �?      �?      �?                      �?      �?      �?              �?                              �?                       @       @              �?       @                       @              �?                      �?                              @      �?              �?                      �?      �?                      4@      l@     �U@      @      E@      @       @      7@                      7@               @                       @      3@      @       @      .@      �?              (@      �?               @                      @      �?               @                       @      �?                      �?               @               @      @              �?                      �?      @              �?                              @                      @      @                      @              @      �?              �?      �?                      �?              �?                      @              0@     �f@      T@      .@      ^@      @@       @      @      @       @      @      @              @      @               @      @               @                              @              �?      @              �?                              @       @              �?                      �?       @                               @              *@     �\@      9@      $@     @\@      9@      $@     �X@      9@      $@     �X@      5@      "@     �G@      ,@      @     �G@      ,@       @     �C@      @              0@      @                      �?              0@      @              "@      @              @      @               @                       @      @                      @               @                      @                      @               @      7@      �?      �?      @                      @              �?                      �?      4@      �?      �?      3@      �?      �?      @                       @              �?      @              �?       @                       @              �?                              �?                      ,@      �?              $@      �?              @                      @      �?                      �?              @                      @                      �?              @       @      "@      @      @       @      �?      @       @      �?      @       @              �?       @                      �?              �?      �?              �?                              �?      �?      @              �?                              @                      @               @                              �?      @                      @              �?       @              �?                               @      @                      �?      J@      @              C@      @               @      @               @       @              @                      �?       @                       @              �?                               @              >@              �?      ,@      @      �?      @      @      �?              @                      @      �?                              @                      $@                              @              ,@              @       @              @                               @              �?     �O@      H@      �?      D@       @              ,@      @              �?      @              �?                              @              *@      �?               @                      @      �?                      �?              @              �?      :@      @              5@      �?              .@                      @      �?              @                      @      �?              @                              �?      �?      @       @                      �?      �?      @      �?      �?       @      �?      �?      �?                      �?              �?                              �?      �?              �?                              �?              @                      7@      D@              "@      @               @      @                      @               @                      @      �?              @                              �?              ,@     �A@              @      :@              @      ,@              @      &@              @      @                      @              @                              @              �?      @                      @              �?                      �?      (@                      (@              �?                      "@      "@              @                      @      "@              @                              "@      @      D@     �a@      @      @@      a@      �?      @      @              @      @               @                      @      @                       @              @      �?              �?      �?              �?                              �?              @              �?              @                       @      �?              �?      �?                                      �?      @      :@     ``@      @      :@     @]@      �?      $@      =@      �?      "@      (@      �?      @      &@              @       @               @                      �?       @                       @              �?              �?      �?      "@      �?               @                      @      �?               @                       @      �?                              �?      �?                      �?              �?                      @      �?              @                              �?              �?      1@              �?      @              �?                              @                      &@      @      0@      V@      @      0@     �U@      @      *@      >@              @      (@              �?      $@              �?       @                      �?              �?      �?              �?                              �?                       @              @       @              @      �?              �?                      @      �?               @      �?                      �?               @                      �?                              �?      @       @      2@              @      @                       @              @      �?              @                      �?      �?                      �?              �?              @      @      .@      @       @      @      @              @                      �?      @              @      @              @                      @      @                                      �?               @                       @      $@              �?       @                       @              �?                      �?       @              �?      @              �?      @                       @              �?      �?              �?                              �?                      @                      �?              @     �L@              �?      C@              �?      @              �?      �?                      �?              �?                              @                      A@               @      3@              �?       @              �?                               @              �?      1@                      *@              �?      @                       @              �?       @              �?                               @       @              �?                      �?       @                                      ,@               @      @              @      �?                      �?              @                      @      @              @                              @      �?     �B@       @      �?      <@      @              6@      @              $@                      (@      @              @                      @      @              @                      @      @                       @              @       @              @                               @      �?      @                      @              �?       @              �?      �?                      �?              �?                              �?                      "@      @                      �?              "@      @              @                      @      @                       @              @      �?               @      �?                      �?               @                       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�BHzhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?       @�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvM�hwh(h+K ��h-��R�(KM���h~�BHW         �                   �`@:��ܕ��?�           ��@       w                    �?V������?�            �u@       R                    �?йS�Ӻ�?�            �n@       5                   �h@��Bkd��?k            `d@                            �?���Q��?0            �Q@                          �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?	       .                   `_@��{d��?-            �P@
       '                    c@໑ɒ��?'             K@       "                    `@`Ӹ����?"            �F@                          �[@4Ea�$t�?             7@                          �Z@�n���?             "@                           �?      �?             @������������������������       �                     �?������������������������       �                     @                          �Z@���Q��?             @������������������������       �                     �?                          `]@      �?             @������������������������       �                     @������������������������       �                     �?                           �?؇���X�?             ,@                           �?ףp=
�?	             $@������������������������       �                     �?                           ]@�����H�?             "@������������������������       �                     @                           I@r�q��?             @                          �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @        !                   `]@      �?             @������������������������       �                     @������������������������       �                     �?#       $                    ^@���7�?             6@������������������������       �                     2@%       &                   `^@      �?             @������������������������       �                     �?������������������������       �                     @(       )                   �U@X�<ݚ�?             "@������������������������       �                      @*       -                   �[@����X�?             @+       ,                   �d@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @/       0                    �?&�q-�?             *@������������������������       �                     @1       4                    `@؇���X�?             @2       3                   @Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @6       ;                    �?�EK	��?;            @W@7       :                   pb@r�q��?             >@8       9                   `t@ ��WV�?             :@������������������������       �                     9@������������������������       �                     �?������������������������       �                     @<       G                   �q@�����?,            �O@=       >                   �[@`Ӹ����?            �F@������������������������       �                     :@?       F                   pk@�KM�]�?             3@@       C                    �?�q�q�?             @A       B                   �]@      �?             @������������������������       �                     �?������������������������       �                     @D       E                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             *@H       I                   �\@�<ݚ�?             2@������������������������       �                      @J       O                    �?      �?             0@K       L                   c@$�q-�?             *@������������������������       �                      @M       N                   �s@z�G�z�?             @������������������������       �                     �?������������������������       �                     @P       Q                   ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @S       `                   @^@��凟��?1            �T@T       U                     �?�h$��W�?             .@������������������������       �                      @V       W                   �W@/y0��k�?             *@������������������������       �                     @X       ]                    �?�n���?             "@Y       \                   @Z@�8��8��?             @Z       [                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @^       _                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @a       p                   �b@��>��M�?)             Q@b       o                    �?0��k���?              J@c       n                   �j@     `�?             @@d       m                    j@     ��?             0@e       l                   @U@hE#߼�?
             .@f       k                    a@�g���e�?             &@g       h                   �]@�8��8��?             @������������������������       �                      @i       j                   P`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �        
             0@������������������������       �                     4@q       r                     �?     ��?	             0@������������������������       �                      @s       v                   @f@X�Cc�?             ,@t       u                   �c@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @x       �                   0i@�H.�!��?<             Y@y       ~                   �[@��/��?            �E@z       }                    �?�g���e�?             &@{       |                   �V@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       �                    �?     0�?             @@������������������������       �                     @�       �                   c@D'�$H{�?             =@�       �                   �_@�*$�Z��?             3@�       �                    @�M�]��?             1@�       �                    �?ƒ_,���?
             .@�       �                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �Q@X�<ݚ�?             "@�       �                    �?      �?              @�       �                   �\@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   `@�z�G��?             $@�       �                    b@�<ݚ�?             "@�       �                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?�P��)�?#            �L@�       �                   P`@.0�w¹�?             E@�       �                   �\@�n���?             B@�       �                   `V@r�q��?             8@������������������������       �                     @�       �                   @\@ԍx�V�?             3@�       �                    Z@r�q��?             2@������������������������       �                     @�       �                     �?      �?             (@������������������������       �                     @�       �                   �`@�q�q�?             "@������������������������       �                      @�       �                   �Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �        	             (@������������������������       �                     @�       �                   @j@��S�ۿ?	             .@�       �                   j@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�                         Pl@6�A��/�?�            @x@�       �                    �?8s�`���?o            `g@�       �                   �c@���;�?,            �Q@�       �                   �_@�N� &�?            �J@�       �                    c@U���N@�?             9@�       �                   �]@Y�����?             6@�       �                   `X@޾�z�<�?             *@�       �                   pa@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    [@ףp=
�?             $@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   h@X�<ݚ�?             "@�       �                    �?z�G�z�?             @�       �                   Pa@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   0a@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?X�Cc�?             <@�       �                   �g@X�<ݚ�?
             2@�       �                    �?�����H�?             "@�       �                   �f@      �?              @�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   @a@�<ݚ�?             "@������������������������       �                     @�       �                    �?�q�q�?             @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �                    �?�ӭ�a��?             2@������������������������       �                     &@�       �                   �d@�$I�$I�?             @������������������������       �                      @�       �                   `f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�c�PFQ�?C             ]@�       �                    _@�h����?             L@�       �                     �?XB���?             =@������������������������       �        	             3@�       �                   �^@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     ;@�                         �c@j�Y�H��?$             N@�       �                    �?��Θ���?"             M@�       �                     �?VUUUUU�?             @������������������������       �                     �?�       �                    k@{�G�z�?             @�       �                    d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �_@8�Z$���?             J@�       �                    _@�t����?	             1@�       �                   �k@z�G�z�?             .@�       �                     �?���!pc�?             &@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @�                          �d@�#-���?            �A@�       �                    b@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     <@������������������������       �                      @      x                  �a@bP�	R��?�             i@      1                   �?�@����?c            @c@                          �?Wj��?&            �L@                        0p@     @�?
             0@������������������������       �                     @      	                  �^@޾�z�<�?             *@������������������������       �                     �?
                        �c@�������?             (@                        �r@�C��2(�?             &@                         �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                        �l@�>$�*��?            �D@������������������������       �                     @      0                  Pe@\�Uo��?             C@                        `a@�!���?             A@������������������������       �                     @                        @[@d��0u��?             >@������������������������       �                      @                         �?��X��?             <@                        �b@؇���X�?             @������������������������       �                     @                        @_@�q�q�?             @������������������������       �                     �?                        �q@      �?              @������������������������       �                     �?������������������������       �                     �?       %                  �[@�ՙ/�?             5@!      "                   �?����X�?             @������������������������       �                     @#      $                  �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @&      -                  �b@և���X�?
             ,@'      (                   ]@�z�G��?             $@������������������������       �                      @)      ,                  @_@      �?              @*      +                  �p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @.      /                   _@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @2      i                  �e@>�HSˏ�?=            @X@3      @                  �m@��r8KP�?4            �U@4      9                   �?8�Z$���?	             *@5      8                   �?�q�q�?             @6      7                  �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?:      ;                  pb@z�G�z�?             $@������������������������       �                     @<      ?                   _@����X�?             @=      >                  0m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @A      b                   @p譎��?+            �R@B      I                   �?<_*{��?'            �P@C      H                  @_@���y4F�?
             3@D      G                  �z@      �?              @E      F                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     &@J      S                    �?�8��8��?             H@K      L                   d@r�q��?             (@������������������������       �                      @M      P                  �d@      �?             @N      O                  p@      �?              @������������������������       �                     �?������������������������       �                     �?Q      R                  @q@      �?              @������������������������       �                     �?������������������������       �                     �?T      a                   �?\��"e��?             B@U      \                   d@t���?             7@V      [                   �?���!pc�?             &@W      Z                  �^@�z�G��?             $@X      Y                  @o@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?]      `                  @_@�8��8��?             (@^      _                  po@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     *@c      h                   �?����X�?             @d      e                  �`@      �?             @������������������������       �                     �?f      g                  �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @j      k                  0n@      �?	             $@������������������������       �                      @l      u                   �?      �?              @m      n                    �?z�G�z�?             @������������������������       �                     �?o      p                   �?      �?             @������������������������       �                     �?q      t                   ]@�q�q�?             @r      s                  pr@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?v      w                  �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @y      �                   �?�R����?            �G@z      �                  �s@�`)j�c�?            �A@{      �                  Pd@8�Z$���?             :@|      �                  �n@��(\���?             4@}      ~                   b@      �?              @������������������������       �                      @      �                  �m@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             (@������������������������       �                     @�      �                  pu@�����H�?             "@�      �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   g@�������?             (@�      �                  hq@�C��2(�?             &@������������������������       �                     "@�      �                  c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�t�b��%      h�h(h+K ��h-��R�(KM�KK��h[�Bh%       �I@     @w@     ps@     �@@      n@     @R@      5@     �g@      A@      0@     @`@      1@      $@      H@      (@               @      �?               @                              �?      $@      G@      &@      "@      D@      @      @      B@      @      @      .@      @      @      @       @      �?      @              �?                              @              @               @                      �?      @              �?      @                                      �?              (@       @              "@      �?              �?                       @      �?              @                      @      �?               @      �?               @                              �?              @                      @      �?              @                              �?              5@      �?              2@                      @      �?                      �?              @              @      @                       @              @       @               @       @                       @               @                      @                      �?      @      @                      @      �?      @              �?       @                       @              �?                              @              @     �T@      @              9@      @              9@      �?              9@                              �?                      @      @     �L@               @     �E@                      :@               @      1@               @      @              �?      @              �?                              @              �?      �?              �?                              �?                      *@              @      ,@               @                       @      ,@              �?      (@                       @              �?      @              �?                              @              �?       @              �?                               @              @     �N@      1@      @      @       @       @                       @      @       @                      @       @      @      @       @      �?      @       @      �?                      �?               @                                      @               @      �?                      �?               @              �?      M@      "@      �?     �G@      @      �?      ;@      @      �?      &@      @      �?      &@      @      �?      @      @      �?       @      @               @              �?              @      �?                                      @              @                      @                              �?              0@                      4@                      &@      @               @                      "@      @              @      @                      @              @                      @              (@     �H@     �C@      &@      ,@      2@      @      �?      @              �?      @              �?                              @      @                      @      *@      .@                      @      @      *@      (@      @      $@      @       @      $@      @       @       @      @       @      @               @                              @                      @      @              @      @               @      @               @                              @              �?                      �?                       @               @                              @      @               @      @               @      �?               @                              �?                      @              �?              �?     �A@      5@      �?      5@      4@      �?      .@      4@      �?      .@       @                      @      �?      .@      @              .@      @              @                      "@      @              @                      @      @                       @              @      �?                      �?              @              �?                                      (@              @                      ,@      �?              @      �?              @                              �?              $@              2@     �`@     �m@      &@      G@     @`@      "@     �@@      =@       @      ?@      ,@       @      *@      @       @      (@       @       @      $@      �?       @      �?                      �?               @                              "@      �?               @      �?                      �?               @                      @              @       @      �?      @              �?       @              �?                      �?       @                       @                       @       @               @                               @                      �?       @              �?                               @              2@      $@               @      $@              �?       @              �?      @              �?      @              �?                              @                      @                      �?              @       @              @                      @       @              �?       @                      �?              �?      �?                      �?              �?                      @                      $@              �?       @      .@                      &@      �?       @      @               @              �?              @                      @      �?                       @      *@     @Y@              �?     �K@              �?      <@                      3@              �?      "@                      "@              �?                              ;@       @      (@      G@       @      $@      G@       @       @       @      �?                      �?       @       @      �?       @              �?                               @                               @               @      F@              @      (@              @      (@              @       @              @                               @                      @               @                      @      @@              @      @              @                              @                      <@               @              @     �U@      [@      @      N@     �V@      �?     �@@      7@      �?      $@      @                      @      �?      $@       @                      �?      �?      $@      �?              $@      �?              @      �?              @                              �?              @              �?                              7@      2@                      @              7@      .@              7@      &@              @                      3@      &@                       @              3@      "@              @      �?              @                       @      �?              �?                      �?      �?                      �?              �?                      *@       @              @       @              @                      �?       @              �?                               @               @      @              @      @                       @              @      �?               @      �?               @                              �?              @                      �?      @              �?                              @                      @       @      ;@      Q@       @      6@     �O@      �?       @      @      �?               @      �?              �?                      �?      �?                                      �?               @       @              @                      @       @              �?       @                       @              �?                      @              �?      ,@     �M@      �?      "@     �L@              @      .@              @      @               @      @                      @               @                       @                              &@      �?      @      E@               @      $@                       @               @       @              �?      �?                      �?              �?                      �?      �?              �?                              �?      �?      @      @@      �?      @      3@              @       @              @      @              @      �?                      �?              @                              @                      �?      �?              &@      �?              @      �?                                      @                      @                      *@              @       @               @       @                      �?               @      �?               @                              �?              @                      @      @               @                      @      @              �?      @                      �?              �?      @                      �?              �?       @              �?      �?                      �?              �?                              �?               @      �?                      �?               @              @      :@      1@      @      0@      0@       @      0@       @       @      0@       @       @      @       @                       @       @      @                      @               @                              (@                              @      �?               @      �?               @                       @      �?                                      @      �?      $@      �?              $@      �?              "@                      �?      �?              �?                              �?      �?                �t�bubhhubehhub.